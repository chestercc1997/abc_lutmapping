module top( V32(0), V32(1), V32(2), V32(3), V56(0), V289(0), V10(0), V13(0), V35(0), V203(0), V288(6), V288(7), V248(0), V249(0), V62(0), V59(0), V174(0), V215(0), V66(0), V70(0), V43(0), V214(0), V37(0), V271(0), V40(0), V45(0), V149(7), V149(6), V149(5), V149(4), V1(0), V7(0), V34(0), V243(0), V244(0), V245(0), V246(0), V247(0), V293(0), V302(0), V270(0), V269(0), V274(0), V202(0), V275(0), V257(7), V257(5), V257(3), V257(1), V257(2), V257(4), V257(6), V9(0), V149(0), V149(1), V149(2), V149(3), V169(1), V165(0), V165(2), V165(4), V165(5), V165(6), V165(7), V165(1), V88(2), V88(3), V55(0), V169(0), V52(0), V5(0), V6(0), V12(0), V11(0), V4(0), V165(3), V51(0), V65(0), V290(0), V279(0), V280(0), V288(4), V288(2), V288(0), V258(0), V229(5), V229(4), V229(3), V229(2), V229(1), V229(0), V223(5), V223(4), V223(3), V223(2), V223(1), V223(0), V189(5), V189(4), V189(3), V189(2), V189(1), V189(0), V183(5), V183(4), V183(3), V183(2), V183(1), V183(0), V239(4), V239(3), V239(2), V239(1), V239(0), V234(4), V234(3), V234(2), V234(1), V234(0), V199(4), V199(3), V199(2), V199(1), V199(0), V194(4), V194(3), V194(2), V194(1), V194(0), V257(0), V32(8), V32(7), V32(6), V32(5), V32(4), V32(11), V32(10), V32(9), V88(1), V88(0), V84(5), V84(4), V84(3), V84(2), V84(1), V84(0), V78(5), V78(4), V2(0), V3(0), V14(0), V213(0), V213(5), V213(4), V213(3), V213(2), V213(1), V268(5), V268(3), V268(1), V268(2), V268(4), V8(0), V60(0), V53(0), V57(0), V109(0), V277(0), V278(0), V259(0), V260(0), V67(0), V68(0), V69(0), V216(0), V175(0), V177(0), V172(0), V171(0), V50(0), V63(0), V71(0), V292(0), V291(0), V91(0), V91(1), V294(0), V207(0), V295(0), V204(0), V205(0), V261(0), V262(0), V100(0), V100(5), V100(4), V100(3), V100(2), V100(1), V240(0), V242(0), V241(0), V33(0), V16(0), V15(0), V101(0), V268(0), V288(1), V288(3), V288(5), V301(0), V108(0), V108(1), V108(2), V108(3), V108(4), V108(5), V124(5), V124(4), V124(3), V124(2), V124(1), V124(0), V132(7), V132(6), V132(5), V132(4), V132(3), V132(2), V132(1), V132(0), V118(5), V118(4), V118(3), V118(2), V118(1), V118(0), V118(7), V118(6), V46(0), V48(0), V102(0), V110(0), V134(1), V134(0), V272(0), V78(2), V78(3), V39(0), V38(0), V42(0), V44(0), V41(0), V78(1), V78(0), V94(0), V94(1), V321(2), V356, V357, V373, V375(0), V377, V393(0), V398(0), V410(0), V423(0), V432, V435(0), V500(0), V508(0), V511(0), V512, V527, V537, V538, V539, V540, V541, V542, V543, V544, V545, V546, V547, V548, V572(9), V572(8), V572(7), V572(6), V572(5), V572(4), V572(3), V572(2), V572(1), V572(0), V585(0), V587, V591(0), V597(0), V603(0), V609(0), V620, V621, V630, V634(0), V640(0), V657, V707, V763, V775, V778, V779, V780, V781, V782, V783, V784, V787, V789, V798(0), V801, V802(0), V821(0), V826(0), V966, V986, V1213(11), V1213(10), V1213(9), V1213(8), V1213(7), V1213(6), V1213(5), V1213(4), V1213(3), V1213(2), V1213(1), V1213(0), V1243(9), V1243(8), V1243(7), V1243(6), V1243(5), V1243(4), V1243(3), V1243(2), V1243(1), V1243(0), V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263, V1264, V1265, V1266, V1267, V1274(0), V1281(0), V1297(4), V1297(3), V1297(2), V1297(1), V1297(0), V1365, V1375, V1378, V1380, V1382, V1384, V1386, V1387, V1392(0), V1423, V1426, V1428, V1429, V1431, V1432, V1439(0), V1440(0), V1451(0), V1459(0), V1467(0), V1470, V1480(0), V1481(0), V1492(0), V1495(0), V1512(3), V1512(2), V1512(1), V1536(0), V1537, V1539, V1552(1), V1552(0), V1613(0), V1613(1), V1620(0), V1629(0), V1645(0), V1652(0), V1669, V1671(0), V1679(0), V1693(0), V1709(4), V1709(3), V1709(2), V1709(1), V1709(0), V1717(0), V1719, V1726(0), V1736, V1741(0), V1745(0), V1757(0), V1758(0), V1759(0), V1760(0), V1771(1), V1771(0), V1781(1), V1781(0), V1829(9), V1829(8), V1829(7), V1829(6), V1829(5), V1829(4), V1829(3), V1829(2), V1829(1), V1829(0), V1832, V1833(0), V1863(0), V1864(0), V1896(0), V1897(0), V1898(0), V1899(0), V1900(0), V1901(0), V1921(5), V1921(4), V1921(3), V1921(2), V1921(1), V1921(0), V1953(1), V1953(7), V1953(6), V1953(5), V1953(4), V1953(3), V1953(2), V1953(0), V1960(1), V1960(0), V1968(0), V1992(1), V1992(0), V650, V651, V652, V653, V654, V655, V656, V1370, V1371, V1372, V1373, V1374 );
  input V32(0), V32(1), V32(2), V32(3), V56(0), V289(0), V10(0), V13(0), V35(0), V203(0), V288(6), V288(7), V248(0), V249(0), V62(0), V59(0), V174(0), V215(0), V66(0), V70(0), V43(0), V214(0), V37(0), V271(0), V40(0), V45(0), V149(7), V149(6), V149(5), V149(4), V1(0), V7(0), V34(0), V243(0), V244(0), V245(0), V246(0), V247(0), V293(0), V302(0), V270(0), V269(0), V274(0), V202(0), V275(0), V257(7), V257(5), V257(3), V257(1), V257(2), V257(4), V257(6), V9(0), V149(0), V149(1), V149(2), V149(3), V169(1), V165(0), V165(2), V165(4), V165(5), V165(6), V165(7), V165(1), V88(2), V88(3), V55(0), V169(0), V52(0), V5(0), V6(0), V12(0), V11(0), V4(0), V165(3), V51(0), V65(0), V290(0), V279(0), V280(0), V288(4), V288(2), V288(0), V258(0), V229(5), V229(4), V229(3), V229(2), V229(1), V229(0), V223(5), V223(4), V223(3), V223(2), V223(1), V223(0), V189(5), V189(4), V189(3), V189(2), V189(1), V189(0), V183(5), V183(4), V183(3), V183(2), V183(1), V183(0), V239(4), V239(3), V239(2), V239(1), V239(0), V234(4), V234(3), V234(2), V234(1), V234(0), V199(4), V199(3), V199(2), V199(1), V199(0), V194(4), V194(3), V194(2), V194(1), V194(0), V257(0), V32(8), V32(7), V32(6), V32(5), V32(4), V32(11), V32(10), V32(9), V88(1), V88(0), V84(5), V84(4), V84(3), V84(2), V84(1), V84(0), V78(5), V78(4), V2(0), V3(0), V14(0), V213(0), V213(5), V213(4), V213(3), V213(2), V213(1), V268(5), V268(3), V268(1), V268(2), V268(4), V8(0), V60(0), V53(0), V57(0), V109(0), V277(0), V278(0), V259(0), V260(0), V67(0), V68(0), V69(0), V216(0), V175(0), V177(0), V172(0), V171(0), V50(0), V63(0), V71(0), V292(0), V291(0), V91(0), V91(1), V294(0), V207(0), V295(0), V204(0), V205(0), V261(0), V262(0), V100(0), V100(5), V100(4), V100(3), V100(2), V100(1), V240(0), V242(0), V241(0), V33(0), V16(0), V15(0), V101(0), V268(0), V288(1), V288(3), V288(5), V301(0), V108(0), V108(1), V108(2), V108(3), V108(4), V108(5), V124(5), V124(4), V124(3), V124(2), V124(1), V124(0), V132(7), V132(6), V132(5), V132(4), V132(3), V132(2), V132(1), V132(0), V118(5), V118(4), V118(3), V118(2), V118(1), V118(0), V118(7), V118(6), V46(0), V48(0), V102(0), V110(0), V134(1), V134(0), V272(0), V78(2), V78(3), V39(0), V38(0), V42(0), V44(0), V41(0), V78(1), V78(0), V94(0), V94(1);
  output V321(2), V356, V357, V373, V375(0), V377, V393(0), V398(0), V410(0), V423(0), V432, V435(0), V500(0), V508(0), V511(0), V512, V527, V537, V538, V539, V540, V541, V542, V543, V544, V545, V546, V547, V548, V572(9), V572(8), V572(7), V572(6), V572(5), V572(4), V572(3), V572(2), V572(1), V572(0), V585(0), V587, V591(0), V597(0), V603(0), V609(0), V620, V621, V630, V634(0), V640(0), V657, V707, V763, V775, V778, V779, V780, V781, V782, V783, V784, V787, V789, V798(0), V801, V802(0), V821(0), V826(0), V966, V986, V1213(11), V1213(10), V1213(9), V1213(8), V1213(7), V1213(6), V1213(5), V1213(4), V1213(3), V1213(2), V1213(1), V1213(0), V1243(9), V1243(8), V1243(7), V1243(6), V1243(5), V1243(4), V1243(3), V1243(2), V1243(1), V1243(0), V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263, V1264, V1265, V1266, V1267, V1274(0), V1281(0), V1297(4), V1297(3), V1297(2), V1297(1), V1297(0), V1365, V1375, V1378, V1380, V1382, V1384, V1386, V1387, V1392(0), V1423, V1426, V1428, V1429, V1431, V1432, V1439(0), V1440(0), V1451(0), V1459(0), V1467(0), V1470, V1480(0), V1481(0), V1492(0), V1495(0), V1512(3), V1512(2), V1512(1), V1536(0), V1537, V1539, V1552(1), V1552(0), V1613(0), V1613(1), V1620(0), V1629(0), V1645(0), V1652(0), V1669, V1671(0), V1679(0), V1693(0), V1709(4), V1709(3), V1709(2), V1709(1), V1709(0), V1717(0), V1719, V1726(0), V1736, V1741(0), V1745(0), V1757(0), V1758(0), V1759(0), V1760(0), V1771(1), V1771(0), V1781(1), V1781(0), V1829(9), V1829(8), V1829(7), V1829(6), V1829(5), V1829(4), V1829(3), V1829(2), V1829(1), V1829(0), V1832, V1833(0), V1863(0), V1864(0), V1896(0), V1897(0), V1898(0), V1899(0), V1900(0), V1901(0), V1921(5), V1921(4), V1921(3), V1921(2), V1921(1), V1921(0), V1953(1), V1953(7), V1953(6), V1953(5), V1953(4), V1953(3), V1953(2), V1953(0), V1960(1), V1960(0), V1968(0), V1992(1), V1992(0), V650, V651, V652, V653, V654, V655, V656, V1370, V1371, V1372, V1373, V1374;
wire n484, n488, n489, n491, n494, n499, n502, n504, n508, n510, n511, n3250, n516, n520, n525, n530, n535, n536, n537, n541, n3412, n549, n550, n554, n555, n556, n557, n558, n559, n587, n595, n597, n599, n609, n611, n3631, n3633, n616, n617, n622, n626, n627, n628, n629, n634, n3832, n647, n651, n652, n658, n661, n667, n668, n675, n678, n681, n694, n701, n707, n710, n716, n720, n725, n739, n745, n746, n752, n758, n764, n773, n781, n789, n792, n797, n801, n806, n811, n816, n820, n825, n832, n834, n839, n843, n848, n852, n4599, n4629, n4631, n856, n866, n871, n878, n4717, n4719, n4720, n4721, n892, n897, n904, n4807, n4809, n4810, n4811, n913, n4874, n4881, n920, n927, n935, n941, n954, n963, n969, n979, n987, n991, n4988, n4994, n4997, n995, n996, n1003, n1011, n1017, n1030, n1039, n1045, n1055, n1063, n1067, n5078, n5084, n5087, n1071, n1073, n1080, n1088, n1094, n1107, n1116, n1122, n1132, n1140, n1144, n5168, n1148, n5214, n5216, n1169, n5339, n5366, n5371, n1173, n1186, n5429, n5451, n5454, n1190, n1203, n5519, n5540, n5544, n1207, n1212, n5586, n5587, n5614, n1218, n1231, n5687, n5726, n1235, n1248, n5816, n1252, n1265, n5878, n1269, n5990, n5992, n1286, n1299, n1304, n1308, n1310, n1311, n1313, n6095, n1318, n1321, n6138, n6223, n1340, n1345, n6359, n1359, n1364, n6495, n1378, n1383, n1389, n6619, n1395, n6693, n1403, n6739, n1409, n6784, n6831, n1421, n1425, n1427, n1430, n6879, n6909, n1451, n7016, n7019, n1456, n1461, n7051, n7053, n1471, n1472, n1474, n7118, n1480, n1489, n1498, n1513, n1522, n1529, n1531, n1532, n1535, n1538, n1539, n1541, n1543, n1546, n7223, n7294, n1566, n1568, n1569, n1573, n1575, n1580, n7378, n7380, n1585, n7475, n7478, n7536, n7539, n7541, n1601, n1605, n1610, n7589, n7618, n1616, n1622, n7640, n1630, n7745, n7746, n1668, n1672, n1679, n1688, n1692, n1702, n1711, n1715, n1725, n8252, n8318, n1746, n1751, n8388, n8454, n1772, n1777, n8524, n8590, n1798, n1803, n1812, n1818, n1824, n1830, n1836, n1842, n1848, n1854, n1856, n1859, n1861, n8946, n1865, n1866, n1868, n1871, n9048, n9087, n9118, n9181, n9228, n1915, n1920, n9304, n9361, n9414, n1949, n1954, n1956, n1964, n9604, n1984, n1989, n1991, n1998, n2007, n9824, n2018, n2024, n2030, n9924, n9953, n2044, n2048, n2054, n10119, n2065, n2071, n2077, n10219, n10248, n2092, n2095, n2101, n10417, n2112, n2118, n2124, n10517, n10546, n2139, n2143, n10663, n10696, n10750, n10941, n2186, n2188, n2212, n11133, n2230, n2231, n2235, n2240, n11355, n2246, n11427, n2249, n2252, n11470, n2254, n11480, n2261, n11541, n2276, n2279, n2282, n11575, n2287, n11605, n11661, n2298, n2307, n2322, n2328, n2338, n11857, n2358, n12005, n2365, n2369, n12134, n12196, n12198, n12263, n12333, n12336, n12337, n12382, n2419, n12414, n12486, n2428, n12496, n2439, n12619, n12703, n12769, n12776, n12818, n2508, n2509, n12891, n12949, n2535, n2571, n2577, n13264, n2587, n13312, n2591, n13382, n13385, n13402, n2605, n13453, n13455, n13513, n13515, n2641, n2647, n2654, n13795, n2670, n2671, n2680, n2689, n2696, n2705, n2714, n2715, n2724, n2733, n2734, n2746, n2755, n2756, n2765, n2774, n2775, n2781, n2789, n2794, n2804, n2811, n2824, n2831, n2834, n2841, n2848, n2851, n15300, n2864, n2868, n2870, n2873, n2880, n15443, n2888, n15455, n15511, n15570, n2904, n2908, n2910, n15681, n15693, n15834, n2960, n2981, n3056, n16040, n16087, n3102, n3103 ; 
assign n484 = (~(n54))*((n55)*((n56)*(n57))) ;
assign n488 = (~(n63))*((~(n61))*((n76)*((n20)*(~(n62))))) ;
assign n489 = (~(n70))*(~(n77)) ;
assign n491 = (~(n54))*((n55)*(~(n56))) ;
assign n494 = ((~(n54))*((n55)*(~(n56))))*((~(n57))*((n27)*(n29))) ;
assign n499 = ((~(n54))*((n55)*(~(n56))))*((~(n57))*((~(n27))*(n29))) ;
assign n502 = (~((n28)*((n30)*((n491)*((~(n57))*((n27)*(n29)))))))*(~((n28)*((n30)*((n491)*((~(n57))*((~(n27))*(n29))))))) ;
assign n504 = (n489)*((~(n68))*(~((~((n28)*((n30)*(n494))))*(~((n28)*((n30)*(n499))))))) ;
assign n508 = (~(n57))*((n56)*((n55)*((n30)*(~(n54))))) ;
assign n510 = (~(n55))*((~(n54))*(~(n56))) ;
assign n511 = (~((~(n57))*((n56)*((n55)*((n30)*(~(n54)))))))*(~((~(n55))*((~(n54))*(~(n56))))) ;
assign n3250 = (((n69)*(~(n183)))*(~(n184)))*(~(n488)) ;
assign n516 = (~((~((n489)*((~(n68))*(~(n502)))))*((~(n508))*(~(n510)))))*(n3250) ;
assign n520 = (n76)*((n62)*((n192)*((n20)*(n64)))) ;
assign n525 = (n60)*((n65)*((n59)*((n63)*((n61)*(n520))))) ;
assign n530 = (n61)*((n76)*((n62)*((n63)*(n64)))) ;
assign n535 = (n60)*((n65)*((n59)*((~(n190))*((n192)*(n530))))) ;
assign n536 = (~(((~((~(n504))*((~(n508))*(~(n510)))))*(n3250))*(n525)))*(~(n535)) ;
assign n537 = (~(n193))*((~(((~((~(n504))*(n511)))*(n3250))*(n525)))*(~(n535))) ;
assign n541 = (~(n57))*((n56)*((n55)*((~(n30))*(~(n54))))) ;
assign n3412 = ((~((~(n57))*((n56)*((n55)*((~(n30))*(~(n54)))))))*(~((~(n54))*((n55)*((n56)*(n57))))))*(~(n5)) ;
assign n549 = (n30)*((n491)*((~(n57))*((n27)*(~(n29))))) ;
assign n550 = (n28)*((n30)*((n491)*((~(n57))*((n27)*(~(n29)))))) ;
assign n554 = (~(n54))*((~(n55))*(n56)) ;
assign n555 = (~((~(n55))*((~(n54))*(~(n56)))))*(~((~(n54))*((~(n55))*(n56)))) ;
assign n556 = (n58)*(~((~((~(n55))*((~(n54))*(~(n56)))))*(~((~(n54))*((~(n55))*(n56)))))) ;
assign n557 = (~(n17))*((~(n55))*((~(n54))*(~(n56)))) ;
assign n558 = (n57)*((~(n17))*((~(n55))*((~(n54))*(~(n56))))) ;
assign n559 = ((n58)*(~((~((~(n55))*((~(n54))*(~(n56)))))*(~((~(n54))*((~(n55))*(n56)))))))*((n57)*((~(n17))*((~(n55))*((~(n54))*(~(n56)))))) ;
assign n587 = (((~((~(n67))*((n66)*(((~(n57))*(n557))*((~(n29))*(~(n30)))))))*(~((n30)*((n29)*((~(n57))*(n557))))))*((~((~(n67))*((n66)*((n29)*((n557)*((~(n30))*(~(n57))))))))*(~((~(n67))*((~(n66))*((n29)*((n557)*((~(n30))*(~(n57))))))))))*(((~((n67)*((n66)*(((~(n57))*(n557))*((~(n29))*(~(n30)))))))*(~((n67)*((~(n66))*((n29)*((n557)*((~(n30))*(~(n57)))))))))*((~((n30)*((~(n29))*((~(n57))*(n557)))))*(~((n67)*((~(n66))*(((~(n57))*(n557))*((~(n29))*(~(n30))))))))) ;
assign n595 = (n57)*((~(n54))*((~(n55))*(n56))) ;
assign n597 = (~(n17))*((~(n57))*((n56)*((n55)*((n30)*(~(n54)))))) ;
assign n599 = (n169)*(~((n168)*((~(n17))*(n508)))) ;
assign n609 = (~((~(n30))*(((~(n54))*((~(n55))*(n56)))*((n29)*(~(n57))))))*((~((n30)*(((~(n54))*((~(n55))*(n56)))*((~(n29))*(~(n57))))))*(~((~(n30))*(((~(n54))*((~(n55))*(n56)))*((~(n29))*(~(n57))))))) ;
assign n611 = (~((n57)*(n557)))*((~((n597)*(~((n169)*(~((n168)*(n597)))))))*(n609)) ;
assign n3631 = ((~((n5)*((n556)*(~(n587)))))*(~((n164)*((n556)*(~(n587))))))*(~(((n587)*(~(n595)))*(n611))) ;
assign n3633 = ((~((~(n166))*((~(n5))*(~(n165)))))*(~((n5)*((n556)*(n558)))))*(~((n164)*((n556)*(n558)))) ;
assign n616 = (~(((n165)*(n537))*(n3412)))*((~(n550))*(~((n3633)*(n3631)))) ;
assign n617 = ((~((~(n504))*(n511)))*(n3250))*((~(n193))*((~(((~((~(n504))*(n511)))*(n3250))*(n525)))*(~(n535)))) ;
assign n622 = (~((~(n57))*((n56)*((n55)*((~(n30))*(~(n54)))))))*(((~((~(n55))*((~(n54))*(~(n56)))))*(~((~(n54))*((~(n55))*(n56)))))*(~((~(n17))*((~(n57))*((n56)*((n55)*((n30)*(~(n54))))))))) ;
assign n626 = ((~((~(n17))*(~(n622))))*(~(((n484)*(~(n599)))*(~((~(n16))*(~(n164)))))))*(~((n484)*(n599))) ;
assign n627 = (~(n16))*((n484)*(~((n169)*(~((n168)*((~(n17))*(n508))))))) ;
assign n628 = (~((~(n54))*((n55)*((n56)*(n57)))))*(~((~(n17))*((~(n57))*((n56)*((n55)*((n30)*(~(n54)))))))) ;
assign n629 = (~((~(n57))*((n56)*((n55)*((~(n30))*(~(n54)))))))*((~((~(n54))*((n55)*((n56)*(n57)))))*(~((~(n17))*((~(n57))*((n56)*((n55)*((n30)*(~(n54))))))))) ;
assign n634 = (~(((~(n541))*(n628))*((n119)*(~((~(n510))*(~(n554)))))))*(~((~((~(n541))*(n628)))*((n129)*((~(n510))*(~(n554)))))) ;
assign n3832 = ((((~(n16))*(n30))*(n484))*(~(n599)))*(n626) ;
assign n647 = (~((~(n626))*((~(n627))*((n537)*(~(n634))))))*((~((n626)*((~(n627))*((n46)*(~(n537))))))*(~((n3832)*(n537)))) ;
assign n651 = (~(n164))*((~(n5))*(~(n16))) ;
assign n652 = ((~((~(n504))*(n511)))*(n3250))*(~((~(n164))*((~(n5))*(~(n16))))) ;
assign n658 = ((n516)*((~(n193))*(n536)))*(((n516)*((~(n193))*(n536)))*(~((~((n3)*((n516)*(~(n651)))))*(~((~((n516)*(~(n651))))*((n134)*(~((n516)*(~(n651)))))))))) ;
assign n661 = (n164)*(~((~((n57)*((~(n54))*((~(n55))*(n56)))))*(~(n597)))) ;
assign n667 = (~(((~((~((~(n617))*((~(n617))*(~(n647)))))*(~(n658))))*(n616))*(~((~(n616))*(~(n661))))))*(~(((n148)*(~(n616)))*((~(n616))*(~(n661))))) ;
assign n668 = (n84)*(n208) ;
assign n675 = (~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))) ;
assign n678 = (~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))) ;
assign n681 = (~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))) ;
assign n694 = (~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))) ;
assign n701 = (~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))) ;
assign n707 = (~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))) ;
assign n710 = (~(((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))))*((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))))*(~((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*(~((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))))) ;
assign n716 = (~(((~(n541))*(n628))*((n95)*(~((~(n510))*(~(n554)))))))*(~((~((~(n541))*(n628)))*((n107)*((~(n510))*(~(n554)))))) ;
assign n720 = (~((n516)*(n537)))*((~(n627))*((n537)*(((~(n617))*(~(n626)))*(~(n716))))) ;
assign n725 = (~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661))))) ;
assign n739 = (n83)*(n209) ;
assign n745 = (n82)*(n210) ;
assign n746 = (~(n11))*(~(n12)) ;
assign n752 = (~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))) ;
assign n758 = (~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))) ;
assign n764 = (~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))) ;
assign n773 = (~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))) ;
assign n781 = (~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))) ;
assign n789 = (~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))) ;
assign n792 = (~((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))))))))))))))*(~(((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758))))))))))*((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))))))))))))) ;
assign n797 = (~(((~(n541))*(n628))*((n97)*(~((~(n510))*(~(n554)))))))*(~((~((~(n541))*(n628)))*((n109)*((~(n510))*(~(n554)))))) ;
assign n801 = (~((n516)*(n537)))*((~(n627))*((n537)*(((~(n617))*(~(n626)))*(~(n797))))) ;
assign n806 = (~((n616)*((~((~(n616))*(~(n661))))*(n801))))*(~(((n1)*(~(n616)))*((~(n616))*(~(n661))))) ;
assign n811 = (~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))) ;
assign n816 = (~(((~(n541))*(n628))*((n96)*(~((~(n510))*(~(n554)))))))*(~((~((~(n541))*(n628)))*((n108)*((~(n510))*(~(n554)))))) ;
assign n820 = (~((n516)*(n537)))*((~(n627))*((n537)*(((~(n617))*(~(n626)))*(~(n816))))) ;
assign n825 = (~((n616)*((~((~(n616))*(~(n661))))*(n820))))*(~(((n2)*(~(n616)))*((~(n616))*(~(n661))))) ;
assign n832 = (~(n30))*((n491)*((n57)*((~(n27))*(~(n29))))) ;
assign n834 = ((~(n70))*(~(n77)))*((~(n28))*(n832)) ;
assign n839 = (~(((~(n541))*(n628))*((n94)*(~((~(n510))*(~(n554)))))))*(~((~((~(n541))*(n628)))*((n106)*((~(n510))*(~(n554)))))) ;
assign n843 = (~((n516)*(n537)))*((~(n627))*((n537)*(((~(n617))*(~(n626)))*(~(n839))))) ;
assign n848 = (~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661))))) ;
assign n852 = (~(n834))*((~((n681)*((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661))))))))*(~((~(n681))*(~((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661)))))))))) ;
assign n4599 = ((n668)*(~((~(n710))*((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661)))))))))*(~((n710)*(~((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661))))))))) ;
assign n4629 = (((((n84)*(n208))*(~((~(n792))*(n806))))*(~((n792)*(~(n806)))))*(~((~(n811))*(n825))))*(~((n811)*(~(n825)))) ;
assign n4631 = ((~((~((~((n681)*(n707)))*(~((~(n681))*(~(n707))))))*(n725)))*(~(((~((n681)*(n707)))*(~((~(n681))*(~(n707)))))*(~(n725)))))*((~(n834))*((~((n681)*(n848)))*(~((~(n681))*(~(n848)))))) ;
assign n856 = (((n4599)*((~((~(n792))*(n806)))*(~((n792)*(~(n806))))))*((~((~(n811))*(n825)))*(~((n811)*(~(n825))))))*(n852) ;
assign n866 = (~((~((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209)))))))))))*(~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))))*(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))) ;
assign n871 = (~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))) ;
assign n878 = (~(n834))*((~((n678)*((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661))))))))*(~((~(n678))*(~((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661)))))))))) ;
assign n4717 = ((n739)*(~(((~((n616)*((~((~(n616))*(~(n661))))*(n801))))*(~(((n1)*(~(n616)))*((~(n616))*(~(n661))))))*(~(n866)))))*(~((~((~((n616)*((~((~(n616))*(~(n661))))*(n801))))*(~(((n1)*(~(n616)))*((~(n616))*(~(n661)))))))*(n866))) ;
assign n4719 = ((n4717)*(~((n825)*(~(n871)))))*(~((~(n825))*(n871))) ;
assign n4720 = (~(((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661))))))*(~((~((n678)*(n701)))*(~((~(n678))*(~(n701))))))))*(~((~((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661)))))))*((~((n678)*(n701)))*(~((~(n678))*(~(n701))))))) ;
assign n4721 = ((~((n725)*(~((~((n678)*(n701)))*(~((~(n678))*(~(n701))))))))*(~((~(n725))*((~((n678)*(n701)))*(~((~(n678))*(~(n701))))))))*((~(n834))*((~((n678)*(n848)))*(~((~(n678))*(~(n848)))))) ;
assign n892 = (~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*(~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))) ;
assign n897 = (~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))) ;
assign n904 = (~(n834))*((~((n675)*((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661))))))))*(~((~(n675))*(~((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661)))))))))) ;
assign n4807 = ((n745)*(~(((~((n616)*((~((~(n616))*(~(n661))))*(n801))))*(~(((n1)*(~(n616)))*((~(n616))*(~(n661))))))*(~(n892)))))*(~((~((~((n616)*((~((~(n616))*(~(n661))))*(n801))))*(~(((n1)*(~(n616)))*((~(n616))*(~(n661)))))))*(n892))) ;
assign n4809 = ((n4807)*(~((n825)*(~(n897)))))*(~((~(n825))*(n897))) ;
assign n4810 = (~(((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661))))))*(~((~((n675)*(n694)))*(~((~(n675))*(~(n694))))))))*(~((~((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661)))))))*((~((n675)*(n694)))*(~((~(n675))*(~(n694))))))) ;
assign n4811 = ((~((n725)*(~((~((n675)*(n694)))*(~((~(n675))*(~(n694))))))))*(~((~(n725))*((~((n675)*(n694)))*(~((~(n675))*(~(n694))))))))*((~(n834))*((~((n675)*(n848)))*(~((~(n675))*(~(n848)))))) ;
assign n913 = (n11)*((n848)*((n806)*((n825)*((~(n725))*(~(n834)))))) ;
assign n4874 = ((~(n746))*(~(n834)))*((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661)))))) ;
assign n4881 = ((((~((~(n11))*(~(n12))))*(n725))*(n806))*(n825))*(n848) ;
assign n920 = (~(n82))*(~(n210)) ;
assign n927 = (~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))) ;
assign n935 = (~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))) ;
assign n941 = (~(((~(n82))*(n210))*(((~(n82))*(n210))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((~(n82))*(n210)))*((~((~(n82))*(n210)))*(~((~(((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))*(~((~((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210)))))))))*(~((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))))))))) ;
assign n954 = (~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~(((~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))) ;
assign n963 = (~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*(~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*(~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(((~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))) ;
assign n969 = (~(((~(n82))*(n210))*(((~(n82))*(n210))*(~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))))))*(~((~((~(n82))*(n210)))*((~((~(n82))*(n210)))*(~((~((~((((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~(((~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))*(~((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*(~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*(~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(((~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))))*(~(((((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~(((~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*(~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*(~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(((~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))))))))) ;
assign n979 = (~(((~(n82))*(n210))*(((~(n82))*(n210))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((~(n82))*(n210)))*((~((~(n82))*(n210)))*(~((~((((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~(((~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))*(~((~(((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))*(~((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~(((~(((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~((~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))))))))) ;
assign n987 = (~(((~(n82))*(n210))*(((~(n82))*(n210))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*(~((~((~(n82))*(n210)))*((~((~(n82))*(n210)))*((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))))))) ;
assign n991 = (~(n834))*((~(((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661))))))*(~(n987))))*(~((~((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661)))))))*(n987)))) ;
assign n4988 = ((~(((~((n616)*((~((~(n616))*(~(n661))))*(n801))))*(~(((n1)*(~(n616)))*((~(n616))*(~(n661))))))*(~(n969))))*(~((~((~((n616)*((~((~(n616))*(~(n661))))*(n801))))*(~(((n1)*(~(n616)))*((~(n616))*(~(n661)))))))*(n969))))*(~(n920)) ;
assign n4994 = ((~((~(n82))*(~(n210))))*(n991))*((~((n725)*(~(n941))))*(~((~(n725))*(n941)))) ;
assign n4997 = (((~((n806)*(~(n969))))*(~((~(n806))*(n969))))*(~((n825)*(~(n979)))))*(~((~(n825))*(n979))) ;
assign n995 = ((((~((n725)*(~(n941))))*(~((~(n725))*(n941))))*(n991))*(n4988))*((~((n825)*(~(n979))))*(~((~(n825))*(n979)))) ;
assign n996 = (~(n83))*(~(n209)) ;
assign n1003 = (~(((n83)*(~(n209)))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((n83)*(~(n209))))))*(~((~((n83)*(~(n209))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((n83)*(~(n209))))))) ;
assign n1011 = (~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*(~((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))))) ;
assign n1017 = (~(((~(n83))*(n209))*(((~(n83))*(n209))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~((~((~(n83))*(n209)))*((~((~(n83))*(n209)))*(~((~(((~(((n83)*(~(n209)))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((n83)*(~(n209))))))*(~((~((n83)*(~(n209))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((n83)*(~(n209))))))))*((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*(~((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))))))))*(~((~((~(((n83)*(~(n209)))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((n83)*(~(n209))))))*(~((~((n83)*(~(n209))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((n83)*(~(n209)))))))))*(~((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*(~((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))))))))))))))) ;
assign n1030 = (~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))*(~(((~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))))) ;
assign n1039 = (~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~((~((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209)))))))))))*(~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))))*(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~(((~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))*(~(((~((~((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209)))))))))))*(~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))))*(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(((~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))))))) ;
assign n1045 = (~(((~(n83))*(n209))*(((~(n83))*(n209))*(~((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))))))))*(~((~((~(n83))*(n209)))*((~((~(n83))*(n209)))*(~((~((~((((~(((n83)*(~(n209)))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((n83)*(~(n209))))))*(~((~((n83)*(~(n209))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((n83)*(~(n209))))))))*((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*(~((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))))))))*((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))*(~(((~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))))))))*(~((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~((~((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209)))))))))))*(~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))))*(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~(((~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))*(~(((~((~((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209)))))))))))*(~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))))*(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(((~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))))))))))*(~(((((~(((n83)*(~(n209)))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((n83)*(~(n209))))))*(~((~((n83)*(~(n209))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((n83)*(~(n209))))))))*((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*(~((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))))))))*((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))*(~(((~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))))))))*((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~((~((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209)))))))))))*(~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))))*(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~(((~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))*(~(((~((~((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209)))))))))))*(~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210)))))))))))*((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))*(~(((~(((~(n11))*(~(n12)))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))*(~((~((~(n11))*(~(n12))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(n11))*(~(n12)))))*((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((n82)*(n210))))))))))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*((~(((n83)*(n209))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((n83)*(n209))))))))))*(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(((~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))))))))))))))) ;
assign n1055 = (~(((~(n83))*(n209))*(((~(n83))*(n209))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))))))*(~((~((~(n83))*(n209)))*((~((~(n83))*(n209)))*(~((~((((~(((n83)*(~(n209)))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((n83)*(~(n209))))))*(~((~((n83)*(~(n209))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((n83)*(~(n209))))))))*((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*(~((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))))))))*((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))*(~(((~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))))))))*(~((~(((~(((n83)*(~(n209)))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((n83)*(~(n209))))))*(~((~((n83)*(~(n209))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((n83)*(~(n209))))))))*((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*(~((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))))))))*(~((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))*(~(((~(((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~(((n83)*(n209))*((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~(((~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))*((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))))))))))))))) ;
assign n1063 = (~(((~(n83))*(n209))*(((~(n83))*(n209))*(~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))*(~((~((~(n83))*(n209)))*((~((~(n83))*(n209)))*((~(((n83)*(~(n209)))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((n83)*(~(n209))))))*(~((~((n83)*(~(n209))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((n83)*(~(n209))))))))))) ;
assign n1067 = (~(n834))*((~(((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661))))))*(~(n1063))))*(~((~((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661)))))))*(n1063)))) ;
assign n5078 = ((~(((~((n616)*((~((~(n616))*(~(n661))))*(n801))))*(~(((n1)*(~(n616)))*((~(n616))*(~(n661))))))*(~(n1045))))*(~((~((~((n616)*((~((~(n616))*(~(n661))))*(n801))))*(~(((n1)*(~(n616)))*((~(n616))*(~(n661)))))))*(n1045))))*(~(n996)) ;
assign n5084 = ((~((~(n83))*(~(n209))))*(n1067))*((~((n725)*(~(n1017))))*(~((~(n725))*(n1017)))) ;
assign n5087 = (((~((n806)*(~(n1045))))*(~((~(n806))*(n1045))))*(~((n825)*(~(n1055)))))*(~((~(n825))*(n1055))) ;
assign n1071 = ((((~((n725)*(~(n1017))))*(~((~(n725))*(n1017))))*(n1067))*(n5078))*((~((n825)*(~(n1055))))*(~((~(n825))*(n1055)))) ;
assign n1073 = (~(n84))*(~(n208)) ;
assign n1080 = (~(((n84)*(~(n208)))*((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*((n84)*(~(n208))))))*(~((~((n84)*(~(n208))))*((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*(~((n84)*(~(n208))))))) ;
assign n1088 = (~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*((~(((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))))*((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))))*(~((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*(~((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))))))))*(~(((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))))*(~((~(((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))))*((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))))*(~((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*(~((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))))))))))))))))))) ;
assign n1094 = (~(((~(n84))*(n208))*(((~(n84))*(n208))*(~((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))))))*(~((~((~(n84))*(n208)))*((~((~(n84))*(n208)))*(~((~(((~(((n84)*(~(n208)))*((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*((n84)*(~(n208))))))*(~((~((n84)*(~(n208))))*((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*(~((n84)*(~(n208))))))))*((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*((~(((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))))*((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))))*(~((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*(~((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))))))))*(~(((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))))*(~((~(((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))))*((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))))*(~((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*(~((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))))))))))))))))))))))*(~((~((~(((n84)*(~(n208)))*((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*((n84)*(~(n208))))))*(~((~((n84)*(~(n208))))*((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*(~((n84)*(~(n208)))))))))*(~((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*((~(((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))))*((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))))*(~((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*(~((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))))))))*(~(((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))))*(~((~(((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))))*((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))))*(~((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*(~((~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694))))))*(~(((~(n83))*(n209))*(~(n675))))))*(~(((~(((n83)*(~(n209)))*(n694)))*(~((~((n83)*(~(n209))))*(~(n694)))))*(((~(n83))*(n209))*(~(n675)))))))))))))))))))))))))))))))))) ;
assign n1107 = (~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758))))))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))))))*(~(((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))))))))))))) ;
assign n1116 = (~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))))))))))))))*(~(((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758))))))))))*((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))))))))*(~(((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))))))))))*(~(((~((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))))))))))))))*(~(((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758))))))))))*((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))))))))))))))*(((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))))))))))) ;
assign n1122 = (~(((~(n84))*(n208))*(((~(n84))*(n208))*(~((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))))))))*(~((~((~(n84))*(n208)))*((~((~(n84))*(n208)))*(~((~((~((((~(((n84)*(~(n208)))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((n84)*(~(n208))))))*(~((~((n84)*(~(n208))))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((n84)*(~(n208))))))))*((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))))*(~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))))))))))))*((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758))))))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))))))*(~(((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))))))))))))))))*(~((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))))))))))))))*(~(((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758))))))))))*((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))))))))*(~(((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))))))))))*(~(((~((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))))))))))))))*(~(((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758))))))))))*((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))))))))))))))*(((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))))))))))))))))))*(~(((((~(((n84)*(~(n208)))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((n84)*(~(n208))))))*(~((~((n84)*(~(n208))))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((n84)*(~(n208))))))))*((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))))*(~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))))))))))))*((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758))))))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))))))*(~(((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))))))))))))*((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))))))))))))))*(~(((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758))))))))))*((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))))))))*(~(((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))))))))))*(~(((~((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))))))))))))))*(~(((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758))))))))))*((~((~(n781))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))))))))*(~((n781)*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*(~(n758))))*((~(((n84)*(n208))*(~(n758))))*(~(((n84)*(n208))*(~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))))))))))))))*(((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))))))))))))))))))) ;
assign n1132 = (~(((~(n84))*(n208))*(((~(n84))*(n208))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*(~((~((~(n84))*(n208)))*((~((~(n84))*(n208)))*(~((~((((~(((n84)*(~(n208)))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((n84)*(~(n208))))))*(~((~((n84)*(~(n208))))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((n84)*(~(n208))))))))*((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))))*(~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))))))))))))*((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758))))))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))))))*(~(((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))))))))))))))))*(~((~(((~(((n84)*(~(n208)))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((n84)*(~(n208))))))*(~((~((n84)*(~(n208))))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((n84)*(~(n208))))))))*((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))))*(~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))))))))))))))))*(~((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758))))))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))))))*(~(((~((((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701)))))))))*((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))*(~((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208))))))))*((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))*(~(((~((((~(n84))*(n208))*(~(n678)))*(~(n701))))*((~(((n84)*(~(n208)))*(~(n701))))*(~((((~(n84))*(n208))*(~(n678)))*((n84)*(~(n208)))))))*(~((~(((n84)*(n208))*(n758)))*(~((~((n84)*(n208)))*(~(n758)))))))))))))*((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*((~(((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678)))))*((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))*(~((~((~(((~(n84))*(n208))*(n678)))*(~((~((~(n84))*(n208)))*(~(n678))))))*(~((~((~(((~(n84))*(n208))*(~(n678))))*(~((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))*(~((((~(n84))*(n208))*(~(n678)))*((~(((n84)*(~(n208)))*(n701)))*(~((~((n84)*(~(n208))))*(~(n701))))))))))))))))))))))))))))) ;
assign n1140 = (~(((~(n84))*(n208))*(((~(n84))*(n208))*(~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))))))))*(~((~((~(n84))*(n208)))*((~((~(n84))*(n208)))*((~(((n84)*(~(n208)))*((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*((n84)*(~(n208))))))*(~((~((n84)*(~(n208))))*((~((~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n675)))*(~((~((~(n83))*(n209)))*(~(n675))))))))))*(~((n84)*(~(n208))))))))))) ;
assign n1144 = (~(n834))*((~(((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661))))))*(~(n1140))))*(~((~((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661)))))))*(n1140)))) ;
assign n5168 = ((~(((~((n616)*((~((~(n616))*(~(n661))))*(n801))))*(~(((n1)*(~(n616)))*((~(n616))*(~(n661))))))*(~(n1122))))*(~((~((~((n616)*((~((~(n616))*(~(n661))))*(n801))))*(~(((n1)*(~(n616)))*((~(n616))*(~(n661)))))))*(n1122))))*(~(n1073)) ;
assign n1148 = ((((~((n725)*(~(n1094))))*(~((~(n725))*(n1094))))*(n1144))*(n5168))*((~((n825)*(~(n1132))))*(~((~(n825))*(n1132)))) ;
assign n5214 = ((((n537)*(~(n834)))*(~(n1148)))*(~((n4629)*(n4631))))*(~((n4881)*(~(n834)))) ;
assign n5216 = ((~((n4719)*(n4721)))*(~((n4809)*(n4811))))*(~((n12)*(n913))) ;
assign n1169 = (~(n834))*((~((~(n681))*((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661))))))))*(~((n681)*(~((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661)))))))))) ;
assign n5339 = ((n668)*(~((~(n707))*((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661)))))))))*(~((n707)*(~((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661))))))))) ;
assign n5366 = ((n84)*(n208))*((~(n834))*((~((~(n681))*(n848)))*(~((n681)*(~(n848)))))) ;
assign n5371 = (((((~((~(n707))*(n725)))*(~((n707)*(~(n725)))))*(~((~(n789))*(n806))))*(~((n789)*(~(n806)))))*(~((~(n764))*(n825))))*(~((n764)*(~(n825)))) ;
assign n1173 = (((n5339)*((~((~(n789))*(n806)))*(~((n789)*(~(n806))))))*(n1169))*((~((~(n764))*(n825)))*(~((n764)*(~(n825))))) ;
assign n1186 = (~(n834))*((~((~(n678))*((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661))))))))*(~((n678)*(~((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661)))))))))) ;
assign n5429 = ((n739)*(~((~(n701))*((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661)))))))))*(~((n701)*(~((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661))))))))) ;
assign n5451 = ((((n83)*(n209))*(~((~(n701))*(n725))))*(~((n701)*(~(n725)))))*(n1186) ;
assign n5454 = (((~((~(n781))*(n806)))*(~((n781)*(~(n806)))))*(~((~(n758))*(n825))))*(~((n758)*(~(n825)))) ;
assign n1190 = (((n5429)*(n1186))*((~((~(n781))*(n806)))*(~((n781)*(~(n806))))))*((~((~(n758))*(n825)))*(~((n758)*(~(n825))))) ;
assign n1203 = (~(n834))*((~((~(n675))*((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661))))))))*(~((n675)*(~((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661)))))))))) ;
assign n5519 = ((n745)*(~((~(n694))*((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661)))))))))*(~((n694)*(~((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661))))))))) ;
assign n5540 = (((n82)*(n210))*(~((~(n773))*(n806))))*(n1203) ;
assign n5544 = ((((~((~(n694))*(n725)))*(~((n694)*(~(n725)))))*(~((n773)*(~(n806)))))*(~((~(n752))*(n825))))*(~((n752)*(~(n825)))) ;
assign n1207 = (((n5519)*(n1203))*((~((~(n773))*(n806)))*(~((n773)*(~(n806))))))*((~((~(n752))*(n825)))*(~((n752)*(~(n825))))) ;
assign n1212 = (n11)*((~(n848))*((~(n725))*((n806)*((n825)*(~(n834)))))) ;
assign n5586 = ((n11)*(n12))*(~((n489)*((~(n28))*(n832)))) ;
assign n5587 = (~((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661)))))))*(n5586) ;
assign n5614 = ((n11)*(~(n834)))*((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661)))))) ;
assign n1218 = (n11)*((n725)*((n806)*((n825)*((~(n834))*(~(n848)))))) ;
assign n1231 = (~(n834))*((~(((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661))))))*(~(n927))))*(~((~((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661)))))))*(n927)))) ;
assign n5687 = ((((~((n725)*(~(n935))))*(~((~(n725))*(n935))))*(~((n806)*(~(n963)))))*(~((~(n806))*(n963))))*((~((n825)*(~(n954))))*(~((~(n825))*(n954)))) ;
assign n5726 = ((n82)*(~(((~((n616)*((~((~(n616))*(~(n661))))*(n801))))*(~(((n1)*(~(n616)))*((~(n616))*(~(n661))))))*(~(n963)))))*(~((~((~((n616)*((~((~(n616))*(~(n661))))*(n801))))*(~(((n1)*(~(n616)))*((~(n616))*(~(n661)))))))*(n963))) ;
assign n1235 = (((n5726)*((~((n725)*(~(n935))))*(~((~(n725))*(n935)))))*(n1231))*((~((n825)*(~(n954))))*(~((~(n825))*(n954)))) ;
assign n1248 = (~(n834))*((~(((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661))))))*(~(n1003))))*(~((~((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661)))))))*(n1003)))) ;
assign n5816 = ((n83)*(~(((~((n616)*((~((~(n616))*(~(n661))))*(n801))))*(~(((n1)*(~(n616)))*((~(n616))*(~(n661))))))*(~(n1039)))))*(~((~((~((n616)*((~((~(n616))*(~(n661))))*(n801))))*(~(((n1)*(~(n616)))*((~(n616))*(~(n661)))))))*(n1039))) ;
assign n1252 = (((n5816)*((~((n725)*(~(n1011))))*(~((~(n725))*(n1011)))))*(n1248))*((~((n825)*(~(n1030))))*(~((~(n825))*(n1030)))) ;
assign n1265 = (~(n834))*((~(((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661))))))*(~(n1080))))*(~((~((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661)))))))*(n1080)))) ;
assign n5878 = (n84)*((~(((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661))))))*(~(n1088))))*(~((~((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661)))))))*(n1088)))) ;
assign n1269 = ((((n5878)*(~((n806)*(~(n1116)))))*(~((~(n806))*(n1116))))*((~((n825)*(~(n1107))))*(~((~(n825))*(n1107)))))*(n1265) ;
assign n5990 = (((n537)*(~(n1269)))*(~((n12)*(n1212))))*(~((n5366)*(n5371))) ;
assign n5992 = ((~((n82)*((n5687)*(n1231))))*(~(n1252)))*(~((n5451)*(n5454))) ;
assign n1286 = (~((n31)*(n53)))*((~((n53)*(n149)))*((~((n32)*(n53)))*(~(((n31)*(n53))*(~((~(n8))*(n167))))))) ;
assign n1299 = (~((n53)*(n150)))*((~((n75)*((n53)*(~((~(n8))*((n44)*(n182)))))))*(~((n53)*(n75)))) ;
assign n1304 = (n60)*((~(n59))*((n10)*(n65))) ;
assign n1308 = (n65)*((n59)*(~(n60))) ;
assign n1310 = (~(n178))*((n200)*(~((n65)*((n59)*(~(n60)))))) ;
assign n1311 = (n120)*(n122) ;
assign n1313 = (n126)*((n124)*((n120)*(n122))) ;
assign n6095 = ((((n121)*(n123))*(n125))*(n127))*(n128) ;
assign n1318 = (n121)*((n123)*((n125)*((n127)*((n128)*(n1313))))) ;
assign n1321 = (n34)*(n35) ;
assign n6138 = ((~(n13))*(n38))*((n37)*((n36)*((n34)*(n35)))) ;
assign n6223 = (~((~((n629)*((n110)*(~((~(n510))*(~(n554)))))))*(~((~(n629))*((n120)*((~(n510))*(~(n554))))))))*(~(n627)) ;
assign n1340 = (~((((~(n626))*(~((n516)*(n537))))*(n537))*(n6223)))*(~(((n136)*((n516)*(n537)))*((n516)*(~(n651))))) ;
assign n1345 = (~((n616)*((~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))*(~(n1340)))))*(~((~(n616))*((n139)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))) ;
assign n6359 = (~((~((n629)*((n112)*(~((~(n510))*(~(n554)))))))*(~((~(n629))*((n122)*((~(n510))*(~(n554))))))))*(~(n627)) ;
assign n1359 = (~((((~(n626))*(~((n516)*(n537))))*(n537))*(n6359)))*(~(((n138)*((n516)*(n537)))*((n516)*(~(n651))))) ;
assign n1364 = (~((n616)*((~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))*(~(n1359)))))*(~((~(n616))*((n141)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))) ;
assign n6495 = (~((~((n629)*((n111)*(~((~(n510))*(~(n554)))))))*(~((~(n629))*((n121)*((~(n510))*(~(n554))))))))*(~(n627)) ;
assign n1378 = (~((((~(n626))*(~((n516)*(n537))))*(n537))*(n6495)))*(~(((n137)*((n516)*(n537)))*((n516)*(~(n651))))) ;
assign n1383 = (~((n616)*((~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))*(~(n1378)))))*(~((~(n616))*((n140)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))) ;
assign n1389 = (n668)*(~(((((n537)*(~(n856)))*(~(n1148)))*(~(n1173)))*(~(n1269)))) ;
assign n6619 = (n537)*(~((((n4807)*(~((n825)*(~(n897)))))*(~((~(n825))*(n897))))*((n4810)*(n904)))) ;
assign n1395 = ((n82)*(n210))*(~((((n6619)*(~(n995)))*(~(n1207)))*(~(n1235)))) ;
assign n6693 = ((~((((n4874)*(n806))*(n825))*(n848)))*(~((((n806)*(n825))*(~(n848)))*(n5587))))*(~((((n5614)*(n806))*(n825))*(~(n848)))) ;
assign n1403 = (n12)*((n11)*(~(((n537)*(~((n12)*(n913))))*(n6693)))) ;
assign n6739 = (n537)*(~((((n4717)*(~((n825)*(~(n871)))))*(~((~(n825))*(n871))))*((n4720)*(n878)))) ;
assign n1409 = ((n83)*(n209))*(~((~(n1190))*(((n6739)*(~(n1071)))*(~(n1252))))) ;
assign n6784 = ((((~(n13))*(n1310))*(~(n1345)))*(~(n1364)))*(~(n1383)) ;
assign n6831 = (~((n6138)*(n1310)))*(~((n1310)*((~(n13))*((n6095)*(n1313))))) ;
assign n1421 = (~(n64))*((n65)*((n59)*(~(n60)))) ;
assign n1425 = (~(n18))*(((~((~(n504))*(n511)))*(n3250))*((n19)*(~(n1308)))) ;
assign n1427 = (n30)*(((~(n54))*((~(n55))*(n56)))*((n29)*(~(n57)))) ;
assign n1430 = (~((n67)*((n66)*((n29)*((n557)*((~(n30))*(~(n57))))))))*(~((~(n67))*((~(n66))*(((~(n57))*(n557))*((~(n29))*(~(n30))))))) ;
assign n6879 = ((~(n17))*(~((n556)*((n57)*((~(n17))*(n510))))))*((~(n1427))*(~((~(n556))*(~(n1430))))) ;
assign n6909 = ((~((n57)*((~(n17))*(n510))))*(n609))*((n587)*(~((n57)*(n554)))) ;
assign n1451 = ((n609)*(~((~((n58)*(~((~(n510))*(~(n554))))))*(~(n587)))))*(~(((n58)*(~((~(n510))*(~(n554)))))*(~(n1430)))) ;
assign n7016 = ((~((~(n489))*(~((n6909)*(n537)))))*(~((n16)*(~((n537)*(n1451))))))*(~((n20)*(~(n537)))) ;
assign n7019 = ((~(n1425))*(~((n5)*(~((n6879)*(~((n556)*(~(n587)))))))))*(~((n15)*((n556)*(~(n587))))) ;
assign n1456 = (((~(n1310))*(~((~(n489))*((~(n599))*(~(n629))))))*(n7016))*(n7019) ;
assign n1461 = (~(n22))*(~((~(n489))*(~((~(n516))*(~((n58)*(~(n555)))))))) ;
assign n7051 = ((((~(n21))*(~((n6138)*(n1310))))*(~((n1304)*(n1310))))*(~((n40)*(n1310))))*(~((n1310)*(n1421))) ;
assign n7053 = ((~((n1310)*((~(n13))*(n1318))))*((~((n1456)*(~((n13)*(n1310)))))*(n1461)))*(n7051) ;
assign n1471 = (n204)*(n205) ;
assign n1472 = (~((~(n204))*(n205)))*(~(n1471)) ;
assign n1474 = (n5)*(~((~(n1427))*(~((~((n58)*(~(n555))))*(~(n1430)))))) ;
assign n7118 = (~((n15)*((n556)*(~(n587)))))*(~((n16)*(~((~((~(n556))*(~(n587))))*((n609)*(~((n556)*(~(n1430))))))))) ;
assign n1480 = (n188)*(~((n5)*(n178))) ;
assign n1489 = (~((~((~((~(n66))*(n67)))*(~((n66)*(~(n67))))))*((~((n139)*(~(n140))))*(~((~(n139))*(n140))))))*(~(((~((~(n66))*(n67)))*(~((n66)*(~(n67)))))*(~((~((n139)*(~(n140))))*(~((~(n139))*(n140))))))) ;
assign n1498 = (~((~((~((n141)*(~(n142))))*(~((~(n141))*(n142)))))*((~((n143)*(~(n144))))*(~((~(n143))*(n144))))))*(~(((~((n141)*(~(n142))))*(~((~(n141))*(n142))))*(~((~((n143)*(~(n144))))*(~((~(n143))*(n144))))))) ;
assign n1513 = (~((~((~((n145)*(~(n146))))*(~((~(n145))*(n146)))))*((~((n147)*(~(n148))))*(~((~(n147))*(n148))))))*(~(((~((n145)*(~(n146))))*(~((~(n145))*(n146))))*(~((~((n147)*(~(n148))))*(~((~(n147))*(n148))))))) ;
assign n1522 = (~((~((~((~(n247))*(n248)))*(~((n247)*(~(n248))))))*((~((n254)*(~(n255))))*(~((~(n254))*(n255))))))*(~(((~((~(n247))*(n248)))*(~((n247)*(~(n248)))))*(~((~((n254)*(~(n255))))*(~((~(n254))*(n255))))))) ;
assign n1529 = (~((~((n257)*((~((~(n1489))*(n1498)))*(~((n1489)*(~(n1498)))))))*(~((~(n257))*(~((~((~(n1489))*(n1498)))*(~((n1489)*(~(n1498))))))))))*(~((~((n256)*((~((~(n1513))*(n1522)))*(~((n1513)*(~(n1522)))))))*(~((~(n256))*(~((~((~(n1513))*(n1522)))*(~((n1513)*(~(n1522)))))))))) ;
assign n1531 = ((~(n54))*((n55)*(~(n56))))*((~(n57))*((~(n27))*(~(n29)))) ;
assign n1532 = (n30)*((n491)*((~(n57))*((~(n27))*(~(n29))))) ;
assign n1535 = (~(n28))*((~(n30))*((n491)*((~(n57))*((n27)*(n29))))) ;
assign n1538 = (n5)*(~((~((n28)*((n30)*(n1531))))*((~((n28)*(n549)))*(~((~(n28))*((~(n30))*(n494))))))) ;
assign n1539 = (~((~(n54))*((~(n55))*(n56))))*(~((~(n17))*((~(n55))*((~(n54))*(~(n56)))))) ;
assign n1541 = (~(n489))*(~((~((~(n17))*(n508)))*((~((~(n54))*((~(n55))*(n56))))*(~((~(n17))*((~(n55))*((~(n54))*(~(n56))))))))) ;
assign n1543 = (~(n1529))*(~((~(n1538))*(~(n1541)))) ;
assign n1546 = (~((n1)*(n789)))*(~((~(n1))*(~(n789)))) ;
assign n7223 = ((((n4)*(~((~(n3))*(~(n707)))))*(~((n3)*(n707))))*(n681))*((~((~(n2))*(~(n764))))*(~((n2)*(n764)))) ;
assign n7294 = ((~((((n3)*((~((n1)*(n789)))*(~((~(n1))*(~(n789))))))*((~((~(n2))*(~(n764))))*(~((n2)*(n764)))))*(n707)))*(~((n764)*((n2)*((~((n1)*(n789)))*(~((~(n1))*(~(n789)))))))))*(~((n1)*(n789))) ;
assign n1566 = (n28)*((~(n30))*((n491)*((~(n57))*((n27)*(n29))))) ;
assign n1568 = (~(n17))*((n28)*((n30)*(n494))) ;
assign n1569 = (~(n30))*((n491)*((~(n57))*((~(n27))*(n29)))) ;
assign n1573 = (n5)*(~(((~((~(n28))*((~(n30))*(n494))))*(~((n28)*((~(n30))*(n494)))))*((~((~(n17))*((n28)*((n30)*(n494)))))*(~((n28)*((~(n30))*(n499))))))) ;
assign n1575 = (~((~(n17))*((~(n55))*((~(n54))*(~(n56))))))*(~((~(n17))*((~(n57))*((n56)*((n55)*((n30)*(~(n54)))))))) ;
assign n1580 = (n28)*((~(n30))*((n491)*((~(n57))*((n27)*(~(n29)))))) ;
assign n7378 = (~((~(n489))*(n554)))*(~((~(n516))*((~(n489))*(~(n1575))))) ;
assign n7380 = ((~((n19)*(n516)))*(~((n19)*(n1580))))*(~(n1573)) ;
assign n1585 = (~((~((n7223)*(n1546)))*(n7294)))*(~((n7380)*(n7378))) ;
assign n7475 = (((~((~(n204))*(n205)))*(~((n204)*(n205))))*(~((n18)*(n19))))*((~(n21))*(~(n22))) ;
assign n7478 = (((~((~(n489))*(~((~(n516))*(~(n556))))))*(n537))*(~(n1543)))*(n7475) ;
assign n7536 = (~((n1310)*((~(n13))*(n1318))))*(((~(n1480))*(~(n1585)))*(n7478)) ;
assign n7539 = (((~((n6138)*(n1310)))*(~((n1304)*(n1310))))*(~((n40)*(n1310))))*(~((n1310)*((~(n64))*(n1308)))) ;
assign n7541 = (n7536)*((n7539)*(~(n1456))) ;
assign n1601 = (~((~(((~(n1389))*(~(n1395)))*((~(n1403))*(~(n1409)))))*(n6784)))*(n7541) ;
assign n1605 = ((n169)*(~((n168)*((~(n17))*(n508)))))*(~((~(n484))*((~(n541))*(~((~(n17))*(n508)))))) ;
assign n1610 = (~(n541))*(~((n202)*(~((~(n484))*(~((~(n17))*(n508))))))) ;
assign n7589 = ((~(n41))*(~((n5)*(n550))))*(~((~(n1610))*((n16)*(n599)))) ;
assign n7618 = (~(n40))*(~((n15)*((n28)*(n549)))) ;
assign n1616 = (~((n7589)*(~((~(n489))*(n1605)))))*(n7618) ;
assign n1622 = (~((n15)*((n28)*((~(n30))*(n494)))))*(~((n5)*(~((~((n28)*((~(n30))*(n494))))*(~((n28)*((~(n30))*(n499)))))))) ;
assign n7640 = (((~((~(n556))*(n558)))*(~((n57)*(n554))))*(~(n484)))*(~(n597)) ;
assign n1630 = (n5)*(~((~((n1535)*(~((~(n1529))*(~((~(n1538))*(~(n1541))))))))*(n7640))) ;
assign n7745 = (((~((n15)*((n556)*(~(n587)))))*(~((n16)*((n556)*(~(n1430))))))*(~((n5)*((~(n556))*(~(n1430))))))*(~((~(n587))*((n16)*(~(n556))))) ;
assign n7746 = (~((n5)*((n30)*((n554)*((n29)*(~(n57)))))))*(~((n16)*(~((~((~(n30))*((n554)*((n29)*(~(n57))))))*((~((n30)*((n554)*((~(n29))*(~(n57))))))*(~((~(n30))*((n554)*((~(n29))*(~(n57))))))))))) ;
assign n1668 = (~(((~(n541))*(n628))*((n93)*(~((~(n510))*(~(n554)))))))*(~((~((~(n541))*(n628)))*((n105)*((~(n510))*(~(n554)))))) ;
assign n1672 = (~((n626)*((~(n627))*((n52)*(~(n537))))))*(~((~(n626))*((~(n627))*((n537)*(~(n1668)))))) ;
assign n1679 = (~((((~((n516)*(n537)))*(~((~(n616))*(~(n661)))))*(n616))*(~(n1672))))*(~(((n135)*(~(n616)))*((~(n616))*(~(n661))))) ;
assign n1688 = (~(((~(n541))*(n628))*((n92)*(~((~(n510))*(~(n554)))))))*(~((~((~(n541))*(n628)))*((n104)*((~(n510))*(~(n554)))))) ;
assign n1692 = (~((n626)*((~(n627))*((n130)*(~(n537))))))*(~((~(n626))*((~(n627))*((n537)*(~(n1688)))))) ;
assign n1702 = (~(((~((~((~(n617))*((~(n617))*(~(n1692)))))*(~((n617)*((n617)*(~(n652)))))))*(n616))*(~((~(n616))*(~(n661))))))*(~(((n134)*(~(n616)))*((~(n616))*(~(n661))))) ;
assign n1711 = (~(((~(n541))*(n628))*((n91)*(~((~(n510))*(~(n554)))))))*(~((~((~(n541))*(n628)))*((n103)*((~(n510))*(~(n554)))))) ;
assign n1715 = (~((n626)*((~(n627))*((n49)*(~(n537))))))*(~((~(n626))*((~(n627))*((n537)*(~(n1711)))))) ;
assign n1725 = (~(((~((~((~(n617))*((~(n617))*(~(n1715)))))*(~((n617)*((n617)*(n652))))))*(n616))*(~((~(n616))*(~(n661))))))*(~(((n133)*(~(n616)))*((~(n616))*(~(n661))))) ;
assign n8252 = ((n50)*(n626))*(~((~(n16))*((n484)*(~(n599))))) ;
assign n8318 = ((~(n626))*(~(n627)))*(~((~((n629)*((n90)*(~(n555)))))*(~((~(n629))*((n102)*(n555)))))) ;
assign n1746 = (~((~((n516)*(n537)))*((~((n516)*(n537)))*(~((~((n8252)*(~(n537))))*(~((n8318)*(n537))))))))*(~(((n516)*(n537))*(((n516)*(n537))*(~((~((n516)*(~(n651))))*(~((~((n516)*(~(n651))))*((n1)*(~((n516)*(~(n651)))))))))))) ;
assign n1751 = (~(((~(n1746))*(n616))*(~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))))*(~((~(n616))*((n132)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))) ;
assign n8388 = ((n48)*(n626))*(~((~(n16))*((n484)*(~(n599))))) ;
assign n8454 = ((~(n626))*(~(n627)))*(~((~((n629)*((n89)*(~(n555)))))*(~((~(n629))*((n101)*(n555)))))) ;
assign n1772 = (~((~((n516)*(n537)))*((~((n516)*(n537)))*(~((~((n8388)*(~(n537))))*(~((n8454)*(n537))))))))*(~(((n516)*(n537))*(((n516)*(n537))*(~((~((n516)*(~(n651))))*(~((~((n516)*(~(n651))))*((n2)*(~((n516)*(~(n651)))))))))))) ;
assign n1777 = (~(((~(n1772))*(n616))*(~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))))*(~((~(n616))*((n131)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))) ;
assign n8524 = ((n51)*(n626))*(~((~(n16))*((n484)*(~(n599))))) ;
assign n8590 = ((~(n626))*(~(n627)))*(~((~((n629)*((n88)*(~(n555)))))*(~((~(n629))*((n100)*(n555)))))) ;
assign n1798 = (~((~((n516)*(n537)))*((~((n516)*(n537)))*(~((~((n8524)*(~(n537))))*(~((n8590)*(n537))))))))*(~(((n516)*(n537))*(((n516)*(n537))*(~((~((n516)*(~(n651))))*(~((~((n516)*(~(n651))))*((n3)*(~((n516)*(~(n651)))))))))))) ;
assign n1803 = (~(((~(n1798))*(n616))*(~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))))*(~((~(n616))*((n138)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))) ;
assign n1812 = (~(((~(n541))*(n628))*((n87)*(~((~(n510))*(~(n554)))))))*(~((~((~(n541))*(n628)))*((n99)*((~(n510))*(~(n554)))))) ;
assign n1818 = (~((n516)*(n537)))*((~((n516)*(n537)))*(~((~((n626)*((~(n627))*((n47)*(~(n537))))))*(~((~(n626))*((~(n627))*((n537)*(~(n1812))))))))) ;
assign n1824 = ((n516)*((~(n193))*(n536)))*(((n516)*((~(n193))*(n536)))*(~((~((n1)*((n516)*(~(n651)))))*(~((~((n516)*(~(n651))))*((n4)*(~((n516)*(~(n651)))))))))) ;
assign n1830 = (~((n616)*((~((~(n616))*(~(n661))))*(~((~(n1818))*(~(n1824)))))))*(~(((n137)*(~(n616)))*((~(n616))*(~(n661))))) ;
assign n1836 = (~(((~(n541))*(n628))*((n86)*(~((~(n510))*(~(n554)))))))*(~((~((~(n541))*(n628)))*((n98)*((~(n510))*(~(n554)))))) ;
assign n1842 = (~((n516)*(n537)))*((~((n516)*(n537)))*(~((~((n626)*((~(n627))*((n52)*(~(n537))))))*(~((~(n626))*((~(n627))*((n537)*(~(n1836))))))))) ;
assign n1848 = ((n516)*((~(n193))*(n536)))*(((n516)*((~(n193))*(n536)))*(~((~((n2)*((n516)*(~(n651)))))*(~((~((n516)*(~(n651))))*((n135)*(~((n516)*(~(n651)))))))))) ;
assign n1854 = (~((n616)*((~((~(n616))*(~(n661))))*(~((~(n1842))*(~(n1848)))))))*(~(((n136)*(~(n616)))*((~(n616))*(~(n661))))) ;
assign n1856 = ((~(n54))*((n55)*((n56)*(n57))))*(~((~(n70))*(~(n77)))) ;
assign n1859 = (n129)*((n6095)*((n126)*((n124)*(n1311)))) ;
assign n1861 = (~(n43))*((n24)*(~((n28)*(n549)))) ;
assign n8946 = ((n244)*(n245))*((n169)*(~((n168)*((~(n17))*(n508))))) ;
assign n1865 = (n244)*((n245)*((n599)*((~(n1859))*(n1861)))) ;
assign n1866 = (~(((~(n599))*(~(n629)))*(n489)))*(~(((n8946)*(~(n1859)))*(n1861))) ;
assign n1868 = ((~(n17))*(n508))*((~((~(n70))*(~(n77))))*(~(n1345))) ;
assign n1871 = (~((~(n70))*(~(n77))))*((~(n17))*(n508)) ;
assign n9048 = ((~((~(n70))*(~(n77))))*(~((n484)*(~(n489)))))*((~(n17))*(n508)) ;
assign n9087 = (~((~((~(n120))*(n121)))*(~((n120)*(~(n121))))))*(~((~((~(n70))*(~(n77))))*((~(n17))*(n508)))) ;
assign n9118 = ((~((~(n70))*(~(n77))))*((~(n17))*(n508)))*(~((n484)*(~(n489)))) ;
assign n9181 = (~((~((n122)*(~((n120)*(n121)))))*(~((~(n122))*((n120)*(n121))))))*(~((~(n489))*((~(n17))*(n508)))) ;
assign n9228 = ((~(n626))*(~(n627)))*(~((~((n629)*((n113)*(~(n555)))))*(~((~(n629))*((n123)*(n555)))))) ;
assign n1915 = (~(((n9228)*(n537))*(~((n516)*(n537)))))*(~(((n516)*(n537))*(((n516)*(n537))*(~((~((n131)*((n516)*(~(n651)))))*(~((~((n516)*(~(n651))))*((n136)*(~((n516)*(~(n651)))))))))))) ;
assign n1920 = (~((n616)*((~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))*(~(n1915)))))*(~((~(n616))*((n142)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))) ;
assign n9304 = ((~((~(n70))*(~(n77))))*(~((n484)*(~(n489)))))*((~(n17))*(n508)) ;
assign n9361 = (~((~((n123)*(~((n121)*((n120)*(n122))))))*(~((~(n123))*((n121)*((n120)*(n122)))))))*(~((~(n489))*(n597))) ;
assign n9414 = ((~(n626))*(~(n627)))*(~((~((n629)*((n114)*(~(n555)))))*(~((~(n629))*((n124)*(n555)))))) ;
assign n1949 = (~(((n9414)*(n537))*(~((n516)*(n537)))))*(~(((n516)*(n537))*(((n516)*(n537))*(~((~((n132)*((n516)*(~(n651)))))*(~((~((n516)*(~(n651))))*((n137)*(~((n516)*(~(n651)))))))))))) ;
assign n1954 = (~((n616)*((~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))*(~(n1949)))))*(~((~(n616))*((n143)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))) ;
assign n1956 = ((~(n17))*(n508))*((~((~(n70))*(~(n77))))*(~(n1954))) ;
assign n1964 = (~(n1856))*(~((~((n124)*(~((n121)*((n123)*((n120)*(n122)))))))*(~((~(n124))*((n121)*((n123)*((n120)*(n122)))))))) ;
assign n9604 = ((~(n626))*(~(n627)))*(~((~((n629)*((n115)*(~(n555)))))*(~((~(n629))*((n125)*(n555)))))) ;
assign n1984 = (~(((n9604)*(n537))*(~((n516)*(n537)))))*(~(((n516)*(n537))*(((n516)*(n537))*(~((~((n133)*((n516)*(~(n651)))))*(~((~((n516)*(~(n651))))*((n138)*(~((n516)*(~(n651)))))))))))) ;
assign n1989 = (~((n616)*((~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))*(~(n1984)))))*(~((~(n616))*((n144)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))) ;
assign n1991 = ((~(n17))*(n508))*((~((~(n70))*(~(n77))))*(~(n1989))) ;
assign n1998 = (~((n125)*(~((n121)*((n123)*((n124)*((n120)*(n122))))))))*(~((~(n125))*((n121)*((n123)*((n124)*((n120)*(n122))))))) ;
assign n2007 = (~(((~(n541))*(n628))*((n116)*(~((~(n510))*(~(n554)))))))*(~((~((~(n541))*(n628)))*((n126)*((~(n510))*(~(n554)))))) ;
assign n9824 = ((((~(n16))*(n27))*(n484))*(~(n599)))*(n626) ;
assign n2018 = (~((n516)*(n537)))*((~((n516)*(n537)))*(~((~((~(n626))*((~(n627))*((n537)*(~(n2007))))))*(~((n9824)*(n537)))))) ;
assign n2024 = ((n516)*((~(n193))*(n536)))*(((n516)*((~(n193))*(n536)))*(~((~((n134)*((n516)*(~(n651)))))*(~((~((n516)*(~(n651))))*((n131)*(~((n516)*(~(n651)))))))))) ;
assign n2030 = (~((n616)*((~((~(n616))*(~(n661))))*(~((~(n2018))*(~(n2024)))))))*(~(((n145)*(~(n616)))*((~(n616))*(~(n661))))) ;
assign n9924 = ((~((~(n70))*(~(n77))))*(~((n484)*(~(n489)))))*((~(n17))*(n508)) ;
assign n9953 = (((~((~(n70))*(~(n77))))*(n27))*(~((~((~(n70))*(~(n77))))*((~(n17))*(n508)))))*(n484) ;
assign n2044 = (~((n126)*(~((n121)*((n123)*((n125)*((n124)*(n1311))))))))*(~((~(n126))*((n121)*((n123)*((n125)*((n124)*(n1311))))))) ;
assign n2048 = (~((n1866)*(n9953)))*(~((~(n1871))*((~(n1866))*((~(n1856))*(~(n2044)))))) ;
assign n2054 = (~(((~(n541))*(n628))*((n117)*(~((~(n510))*(~(n554)))))))*(~((~((~(n541))*(n628)))*((n127)*((~(n510))*(~(n554)))))) ;
assign n10119 = ((((~(n16))*(n28))*(n484))*(~(n599)))*(n626) ;
assign n2065 = (~((n516)*(n537)))*((~((n516)*(n537)))*(~((~((~(n626))*((~(n627))*((n537)*(~(n2054))))))*(~((n10119)*(n537)))))) ;
assign n2071 = ((n516)*((~(n193))*(n536)))*(((n516)*((~(n193))*(n536)))*(~((~((n135)*((n516)*(~(n651)))))*(~((~((n516)*(~(n651))))*((n132)*(~((n516)*(~(n651)))))))))) ;
assign n2077 = (~((n616)*((~((~(n616))*(~(n661))))*(~((~(n2065))*(~(n2071)))))))*(~(((n146)*(~(n616)))*((~(n616))*(~(n661))))) ;
assign n10219 = ((~((~(n70))*(~(n77))))*(~((n484)*(~(n489)))))*((~(n17))*(n508)) ;
assign n10248 = (((~((~(n70))*(~(n77))))*(n28))*(~((~((~(n70))*(~(n77))))*((~(n17))*(n508)))))*(n484) ;
assign n2092 = (~(n1856))*(~((~((n127)*(~((n121)*((n123)*((n125)*(n1313)))))))*(~((~(n127))*((n121)*((n123)*((n125)*(n1313)))))))) ;
assign n2095 = (~((n1866)*(n10248)))*(~((~(n1871))*((~(n1866))*(n2092)))) ;
assign n2101 = (~(((~(n541))*(n628))*((n118)*(~((~(n510))*(~(n554)))))))*(~((~((~(n541))*(n628)))*((n128)*((~(n510))*(~(n554)))))) ;
assign n10417 = ((((~(n16))*(n29))*(n484))*(~(n599)))*(n626) ;
assign n2112 = (~((n516)*(n537)))*((~((n516)*(n537)))*(~((~((~(n626))*((~(n627))*((n537)*(~(n2101))))))*(~((n10417)*(n537)))))) ;
assign n2118 = ((n516)*((~(n193))*(n536)))*(((n516)*((~(n193))*(n536)))*(~((~((n4)*((n516)*(~(n651)))))*(~((~((n516)*(~(n651))))*((n133)*(~((n516)*(~(n651)))))))))) ;
assign n2124 = (~((n616)*((~((~(n616))*(~(n661))))*(~((~(n2112))*(~(n2118)))))))*(~(((n147)*(~(n616)))*((~(n616))*(~(n661))))) ;
assign n10517 = ((~((~(n70))*(~(n77))))*(~((n484)*(~(n489)))))*((~(n17))*(n508)) ;
assign n10546 = (((~((~(n70))*(~(n77))))*(n29))*(~((~((~(n70))*(~(n77))))*((~(n17))*(n508)))))*(n484) ;
assign n2139 = (~((n128)*(~((n121)*((n123)*((n125)*((n127)*(n1313))))))))*(~((~(n128))*((n121)*((n123)*((n125)*((n127)*(n1313))))))) ;
assign n2143 = (~((n1866)*(n10546)))*(~((~(n1871))*((~(n1866))*((~(n1856))*(~(n2139)))))) ;
assign n10663 = ((~((~(n70))*(~(n77))))*(~((n484)*(~(n489)))))*((~(n17))*(n508)) ;
assign n10696 = (((~((~(n70))*(~(n77))))*(n30))*(~((~((~(n70))*(~(n77))))*((~(n17))*(n508)))))*(n484) ;
assign n10750 = ((~((n484)*(~(n489))))*(~((~(n489))*(n597))))*(~((~((n129)*(~((n6095)*(n1313)))))*(~((~(n129))*((n6095)*(n1313)))))) ;
assign n10941 = ((~((n65)*((n59)*(~(n60)))))*(n16))*(~(n22)) ;
assign n2186 = (~((~(n559))*(~((n1535)*(~((~(n1529))*(~((~(n1538))*(~(n1541))))))))))*(n10941) ;
assign n2188 = ((n28)*((~(n30))*(n494)))*((n15)*(~(n22))) ;
assign n2212 = (n246)*(((~(n70))*(~(n77)))*((n201)*((n244)*(n245)))) ;
assign n11133 = (((n201)*(~((~(n541))*((~(n484))*(~(n597))))))*(~((n5)*(~((~(n484))*(~(n597)))))))*(n489) ;
assign n2230 = (n18)*((n172)*(n178)) ;
assign n2231 = (~(n28))*((~(n30))*((n491)*((~(n57))*((~(n27))*(n29))))) ;
assign n2235 = (~(n556))*((~((~(n28))*(n1569)))*((~(n1568))*((~(n554))*(n1480)))) ;
assign n2240 = (n15)*((n1480)*((~(n554))*((~(n28))*((~(n30))*(n499))))) ;
assign n11355 = ((~((n16)*((n1480)*((~(n554))*(n556)))))*(~((~(n556))*((~(n2231))*((~(n1568))*((~(n554))*(n1480)))))))*(~(((n16)*(n1568))*((~(n554))*(n1480)))) ;
assign n2246 = (~(n2240))*(((~(n2230))*(~(n22)))*(n11355)) ;
assign n11427 = (~((n489)*((~(n1610))*((n192)*(~(n599))))))*(~((n599)*((~(n45))*((n246)*((n489)*((n192)*(~(n1610)))))))) ;
assign n2249 = (~((n11133)*(~(n599))))*((n2246)*((n11427)*(~((n599)*((~(n45))*(n2212)))))) ;
assign n2252 = (n64)*((~(n79))*((n65)*((n59)*(~(n60))))) ;
assign n11470 = (~((n64)*((~(n79))*((n65)*((n59)*(~(n60)))))))*(~(n1421)) ;
assign n2254 = (n2249)*((n11470)*(~(n40))) ;
assign n11480 = ((n20)*(n151))*(~(n536)) ;
assign n2261 = (n5)*(~((~((n28)*((n30)*(n494))))*(~((n28)*((n30)*(n499)))))) ;
assign n11541 = (~((~(n1308))*((n16)*((n1480)*((~(n554))*(n556))))))*(~((~(n1308))*(((n16)*(n1568))*((~(n554))*(n1480))))) ;
assign n2276 = ((~((n79)*(n1308)))*(~(n2240)))*((n11541)*(~((~(n1308))*(n2235)))) ;
assign n2279 = (~(n28))*((~(n30))*((n491)*((~(n57))*((n27)*(~(n29)))))) ;
assign n2282 = (n28)*((~(n30))*((n491)*((~(n57))*((~(n27))*(~(n29)))))) ;
assign n11575 = (((~(n16))*(n85))*(~(n170)))*(~(n171)) ;
assign n2287 = (~(n28))*((n30)*((n491)*((~(n57))*((~(n27))*(~(n29)))))) ;
assign n11605 = (((((~((n28)*((n30)*((n491)*((~(n57))*((~(n27))*(~(n29))))))))*(~((~(n28))*((~(n30))*((n491)*((~(n57))*((n27)*(~(n29)))))))))*(~((~(n28))*((n30)*((n491)*((~(n57))*((n27)*(~(n29)))))))))*(~((n28)*((~(n30))*((n491)*((~(n57))*((~(n27))*(~(n29)))))))))*(~((~(n28))*((n30)*((n491)*((~(n57))*((~(n27))*(~(n29)))))))))*(~((~(n28))*((n30)*((n491)*((~(n57))*((n27)*(n29))))))) ;
assign n11661 = (~((n15)*(~((~((~(n28))*((~(n30))*(n494))))*(~((n28)*((~(n30))*(n499))))))))*(~((n78)*((n28)*((~(n30))*(n494))))) ;
assign n2298 = (~((n5)*(~((~((~((~(n193))*(n536)))*(n11575)))*(n11605)))))*(n11661) ;
assign n2307 = (~(n22))*(~((~((~(n541))*(~((n202)*(~(n628))))))*(~((~(n1304))*(n2254))))) ;
assign n2322 = (~(n28))*((~(n30))*((n491)*((n57)*((n27)*(~(n29)))))) ;
assign n2328 = (~((~(n28))*((~(n30))*((n491)*((~(n57))*((~(n27))*(~(n29))))))))*((~((~(n28))*((n29)*((n491)*((n30)*((~(n27))*(~(n57))))))))*(~((~((n28)*((~(n30))*((n491)*((n57)*((~(n27))*(~(n29))))))))*((n57)*((n491)*((~((~(n28))*((~(n30))*((n491)*((n57)*((~(n27))*(~(n29))))))))*(~((~(n28))*((~(n30))*((n491)*((n57)*((n27)*(~(n29)))))))))))))) ;
assign n2338 = (~((~((n55)*((n54)*(~(n56)))))*((n2328)*((~((n55)*((n54)*(n56))))*(~((n56)*((n54)*(~(n55)))))))))*((n537)*(~((~(n40))*(~(n2328))))) ;
assign n11857 = ((((~(n6))*(~(n40)))*(n151))*(~((n64)*((~(n79))*(n1308)))))*(~((n79)*(~(n1308)))) ;
assign n2358 = (~((~(n70))*(~((~(n17))*((n5)*(~(n502)))))))*((~(n502))*((n5)*(n516))) ;
assign n12005 = ((~((n5)*(~(n2328))))*(~((n488)*(~(n502)))))*(~(n2358)) ;
assign n2365 = (n16)*(~(((~((~(n556))*(n558)))*(~(n595)))*(n629))) ;
assign n2369 = (~(n2358))*(((~((~(n537))*(n11575)))*(n11605))*((n5)*(n2328))) ;
assign n12134 = (((~((n57)*((~(n17))*(n510))))*(~((n57)*(n554))))*(~(n597)))*(n609) ;
assign n12196 = ((~(n9))*(~(n17)))*(n73) ;
assign n12198 = ((n12196)*(n149))*(~(((n28)*(n549))*(~((~(n164))*(~(n181)))))) ;
assign n12263 = ((~(n1427))*(~((~(n556))*(n558))))*(~(n484)) ;
assign n12333 = ((n16)*(~(n1310)))*(((~(n541))*(~(n595)))*(~((~(n556))*(~(n1430))))) ;
assign n12336 = ((~((~(n17))*((n28)*((n30)*(n494)))))*(~((~(n28))*(n832))))*(~((~(n17))*((n28)*((n30)*(n499))))) ;
assign n12337 = (n12336)*((n151)*((n12263)*(~(n597)))) ;
assign n12382 = (~(((n58)*(~((~((~(n55))*((~(n54))*(~(n56)))))*(~((~(n54))*((~(n55))*(n56)))))))*((~(n17))*((~(n55))*((~(n54))*(~(n56)))))))*(~((~(n40))*((~(n54))*((~(n55))*(n56))))) ;
assign n2419 = ((n12382)*(~((~(n17))*((n28)*((n30)*(n494))))))*(~((~(n28))*((~(n30))*(n499)))) ;
assign n12414 = (((~(n6))*(n151))*((n188)*(~((n5)*(n178)))))*(~(n1308)) ;
assign n12486 = (((~((n28)*((n30)*(n499))))*(~(n1308)))*(n508))*(n1480) ;
assign n2428 = (n508)*((n79)*((n65)*((n59)*(~(n60))))) ;
assign n12496 = (n152)*((n151)*(~((n5)*(n2279)))) ;
assign n2439 = (~(n1480))*(~((~(n63))*((~(n61))*((~(n76))*((~(n62))*(~(n64))))))) ;
assign n12619 = ((((n15)*(n609))*(~((~(n556))*(~(n587)))))*(~((n556)*(~(n1430)))))*(n537) ;
assign n12703 = (((~(n1859))*(~((n13)*(n489))))*(n489))*(n541) ;
assign n12769 = ((~((n13)*(n489)))*(~(n628)))*(~((n489)*(n1859))) ;
assign n12776 = (~(((~((n489)*((~(n1610))*((n192)*(~(n599))))))*(~(n599)))*(n12703)))*(~((~((n489)*((~(n1610))*((n192)*(~(n599))))))*((n12769)*(~((n489)*(n599)))))) ;
assign n12818 = (((n5)*(n32))*((n28)*(n1532)))*(~(n1308)) ;
assign n2508 = (~(n15))*((~(n5))*(~(n180))) ;
assign n2509 = (~((~(n193))*(n536)))*(~((~(n15))*((~(n5))*(~(n180))))) ;
assign n12891 = ((((n20)*(~(n61)))*(~(n62)))*(n63))*(n76) ;
assign n12949 = ((n78)*(~((n28)*((~(n30))*(n494)))))*(~((n556)*(~(n587)))) ;
assign n2535 = (n207)*((n162)*((n161)*((n160)*((n158)*(n159))))) ;
assign n2571 = (~((~(n174))*((~(n19))*((~(n20))*(~(n173))))))*((n18)*(n151)) ;
assign n2577 = (~(((~(n54))*((~(n55))*(n56)))*(n1480)))*(~((n27)*((n5)*((~(n54))*((~(n55))*(n56)))))) ;
assign n13264 = (((~((n5)*(n178)))*(~(n13)))*(n177))*(~((n179)*((n5)*(~(n555))))) ;
assign n2587 = (~((n16)*((n556)*(~(n1430)))))*(~((~((n169)*(~(n629))))*(n13264))) ;
assign n13312 = (n2577)*(~((~((~(n178))*(n1474)))*((~((~(n24))*(~(n43))))*(n2587)))) ;
assign n2591 = (n13312)*(n2249) ;
assign n13382 = ((~((n4629)*(n4631)))*(~((n4719)*(n4721))))*(~((n4809)*(n4811))) ;
assign n13385 = (((~((n12)*(n913)))*(~(n1190)))*(~((n12)*(n1212))))*(~((n5366)*(n5371))) ;
assign n13402 = (~(n2261))*(~((~((n554)*(n1480)))*(~((n27)*((n5)*(n554)))))) ;
assign n2605 = (~((n5366)*(n5371)))*(~(n1269)) ;
assign n13453 = ((~((n4629)*(n4631)))*(~((n4809)*(n4811))))*(~((n4994)*(n4997))) ;
assign n13455 = ((~(n1148))*(~((n5540)*(n5544))))*(~((n82)*((n5687)*(n1231)))) ;
assign n13513 = ((~((n4629)*(n4631)))*(~((n4719)*(n4721))))*(~((n5084)*(n5087))) ;
assign n13515 = ((~(n1148))*(~((n5451)*(n5454))))*(~(n1252)) ;
assign n2641 = (((~((~((n110)*(~(n111))))*(~((~(n110))*(n111)))))*(~((~(n489))*(~(n1539)))))*(n595))*(n489) ;
assign n2647 = (~((n28)*(n832)))*((~((~(n28))*(n549)))*((n230)*((~(n28))*(n1532)))) ;
assign n2654 = (~((~((n28)*(n832)))*((~((~(n28))*(n549)))*((n231)*((~(n28))*(n1532))))))*(~(((n28)*(n832))*((~((~(n28))*(n549)))*((n217)*(~((~(n28))*(n1532))))))) ;
assign n13795 = (~((~(n28))*((~(n30))*((n491)*((~(n57))*((n27)*(~(n29))))))))*((~((n28)*((~(n30))*((n491)*((~(n57))*((~(n27))*(~(n29))))))))*(~((~(n28))*((~(n30))*((n491)*((n57)*((n27)*(~(n29))))))))) ;
assign n2670 = (~((~(n2322))*((~(n2287))*((~(n2279))*((n195)*(n2282))))))*(~((~(n2322))*((~(n2287))*((n2279)*((n153)*(~(n2282))))))) ;
assign n2671 = (~((n218)*((n13795)*(n2287))))*(n2670) ;
assign n2680 = (~((~(n2322))*((n2287)*((~(n2279))*((n219)*(~(n2282)))))))*(~((n2322)*((~(n2287))*((~(n2279))*((n216)*(~(n2282))))))) ;
assign n2689 = (~((~(n2322))*((~(n2287))*((~(n2279))*((n196)*(n2282))))))*(~((~(n2322))*((~(n2287))*((n2279)*((n154)*(~(n2282))))))) ;
assign n2696 = (~((~((~((n2647)*(n2654)))*(~((~(n2647))*(~(n2654))))))*((~((~(n2671))*((n2680)*(n2689))))*(~((n2671)*(~((n2680)*(n2689))))))))*(~(((~((n2647)*(n2654)))*(~((~(n2647))*(~(n2654)))))*(~((~((~(n2671))*((n2680)*(n2689))))*(~((n2671)*(~((n2680)*(n2689))))))))) ;
assign n2705 = (~((~(n2322))*((n2287)*((~(n2279))*((n220)*(~(n2282)))))))*(~((n2322)*((~(n2287))*((~(n2279))*((n215)*(~(n2282))))))) ;
assign n2714 = (~((~(n2322))*((~(n2287))*((~(n2279))*((n197)*(n2282))))))*(~((~(n2322))*((~(n2287))*((n2279)*((n155)*(~(n2282))))))) ;
assign n2715 = (n2705)*(n2714) ;
assign n2724 = (~((~(n2322))*((n2287)*((~(n2279))*((n221)*(~(n2282)))))))*(~((n2322)*((~(n2287))*((~(n2279))*((n214)*(~(n2282))))))) ;
assign n2733 = (~((~(n2322))*((~(n2287))*((~(n2279))*((n198)*(n2282))))))*(~((~(n2322))*((~(n2287))*((n2279)*((n156)*(~(n2282))))))) ;
assign n2734 = (n2724)*(n2733) ;
assign n2746 = (~((~(n2322))*((n2287)*((~(n2279))*((n222)*(~(n2282)))))))*(~((n2322)*((~(n2287))*((~(n2279))*((n213)*(~(n2282))))))) ;
assign n2755 = (~((~(n2322))*((~(n2287))*((~(n2279))*((n199)*(n2282))))))*(~((~(n2322))*((~(n2287))*((n2279)*((n157)*(~(n2282))))))) ;
assign n2756 = (n2746)*(n2755) ;
assign n2765 = (~((~(n2322))*((n2287)*((~(n2279))*((n223)*(~(n2282)))))))*(~((n2322)*((~(n2287))*((~(n2279))*((n212)*(~(n2282))))))) ;
assign n2774 = (~((~(n2322))*((~(n2287))*((~(n2279))*((n194)*(n2282))))))*(~((~(n2322))*((~(n2287))*((n2279)*((n152)*(~(n2282))))))) ;
assign n2775 = (n2765)*(n2774) ;
assign n2781 = (~((~((~((~(n2715))*(n2734)))*(~((n2715)*(~(n2734))))))*((~((~(n2756))*(n2775)))*(~((n2756)*(~(n2775)))))))*(~(((~((~(n2715))*(n2734)))*(~((n2715)*(~(n2734)))))*(~((~((~(n2756))*(n2775)))*(~((n2756)*(~(n2775)))))))) ;
assign n2789 = (~((n238)*(((~(n1566))*(~((n28)*(n1569))))*((~(n28))*(n549)))))*(~((n240)*((~((~(n1566))*(~((n28)*(n1569)))))*(~((~(n28))*(n549)))))) ;
assign n2794 = (~((n239)*(((~(n1566))*(~((n28)*(n1569))))*((~(n28))*(n549)))))*(~((n241)*((~((~(n1566))*(~((n28)*(n1569)))))*(~((~(n28))*(n549)))))) ;
assign n2804 = (~((~((n28)*(n832)))*((~((~(n28))*(n549)))*((n224)*((~(n28))*(n1532))))))*(~((~((n28)*(n832)))*(((~(n28))*(n549))*((n232)*(~((~(n28))*(n1532))))))) ;
assign n2811 = (~((~((n28)*(n832)))*((~((~(n28))*(n549)))*((n225)*((~(n28))*(n1532))))))*(~((~((n28)*(n832)))*(((~(n28))*(n549))*((n233)*(~((~(n28))*(n1532))))))) ;
assign n2824 = (~((~((n28)*(n832)))*((~((~(n28))*(n549)))*((n226)*((~(n28))*(n1532))))))*(~((~((n28)*(n832)))*(((~(n28))*(n549))*((n234)*(~((~(n28))*(n1532))))))) ;
assign n2831 = (~((~((n28)*(n832)))*((~((~(n28))*(n549)))*((n227)*((~(n28))*(n1532))))))*(~((~((n28)*(n832)))*(((~(n28))*(n549))*((n235)*(~((~(n28))*(n1532))))))) ;
assign n2834 = (~((~(n2824))*(n2831)))*(~((n2824)*(~(n2831)))) ;
assign n2841 = (~((~((n28)*(n832)))*((~((~(n28))*(n549)))*((n228)*((~(n28))*(n1532))))))*(~((~((n28)*(n832)))*(((~(n28))*(n549))*((n236)*(~((~(n28))*(n1532))))))) ;
assign n2848 = (~((~((n28)*(n832)))*((~((~(n28))*(n549)))*((n229)*((~(n28))*(n1532))))))*(~((~((n28)*(n832)))*(((~(n28))*(n549))*((n237)*(~((~(n28))*(n1532))))))) ;
assign n2851 = (~((~(n2841))*(n2848)))*(~((n2841)*(~(n2848)))) ;
assign n15300 = (~((n17)*((n65)*((n59)*(~(n60))))))*(~((~(n40))*(n183))) ;
assign n2864 = (~(n187))*(~((n28)*((~(n30))*(n494)))) ;
assign n2868 = (~((n15)*(n186)))*(~((n16)*(n185))) ;
assign n2870 = ((~((~(n26))*(n253)))*(~((n26)*(~(n253)))))*(~((n1535)*(~(n2868)))) ;
assign n2873 = (~((n12414)*(~(n2419))))*(~((n27)*((~((~(n70))*(~(n77))))*(n554)))) ;
assign n2880 = (~(n6))*((~(n64))*((n65)*((n59)*(~(n60))))) ;
assign n15443 = (~((n85)*((~(n171))*((~(n16))*(~(n170))))))*(n151) ;
assign n2888 = (n536)*(~((n193)*((n15443)*(n193)))) ;
assign n15455 = (((((~((n28)*((n30)*((n491)*((~(n57))*((~(n27))*(~(n29))))))))*(~((~(n28))*((~(n30))*((n491)*((~(n57))*((n27)*(~(n29)))))))))*(~((~(n28))*((n30)*((n491)*((~(n57))*((n27)*(~(n29)))))))))*(~((n28)*((~(n30))*((n491)*((~(n57))*((~(n27))*(~(n29)))))))))*(~((~(n28))*((n30)*((n491)*((~(n57))*((~(n27))*(~(n29)))))))))*(~((~(n28))*((n30)*((n491)*((~(n57))*((n27)*(n29))))))) ;
assign n15511 = (~((n28)*((~(n30))*((n491)*((~(n57))*((n27)*(n29)))))))*((~((~(n28))*((~(n30))*((n491)*((~(n57))*((n27)*(n29)))))))*(~((n28)*((~(n30))*((n491)*((~(n57))*((~(n27))*(n29)))))))) ;
assign n15570 = ((~(n6))*(~(n2252)))*(~(((n15511)*((n15455)*(n2888)))*(n2888))) ;
assign n2904 = (~((n19)*(n1580)))*(~((~(n6))*((~(n2276))*((n15455)*(n2888))))) ;
assign n2908 = (~((~(n54))*((n55)*(~(n56)))))*(~((~(n55))*((~(n54))*(~(n56))))) ;
assign n2910 = (n79)*((n1308)*(~((~((~(n54))*((n55)*(~(n56)))))*(~((~(n55))*((~(n54))*(~(n56)))))))) ;
assign n15681 = (((~(n2908))*(~(n1308)))*(n1480))*(~((n28)*((n30)*(n499)))) ;
assign n15693 = (n194)*((n151)*(~((n5)*(n2282)))) ;
assign n15834 = ((((~(n178))*(n200))*(~((~(n81))*(n595))))*(~(n1304)))*(~(n1308)) ;
assign n2960 = (~((n57)*(n554)))*(~((~((n169)*(~((n168)*(n597)))))*(~(n629)))) ;
assign n2981 = (~((n508)*((n204)*(~(n205)))))*(~(((~(n55))*((~(n54))*(~(n56))))*((n204)*(~(n205))))) ;
assign n3056 = (n5)*(n2322) ;
assign n16040 = ((~((n206)*((~(n216))*((~(n204))*(n205)))))*(n151))*(n243) ;
assign n16087 = ((~(n55))*((~(n54))*(~(n56))))*(~((~(n242))*((~((~(n204))*(n205)))*(~((n204)*(~(n205))))))) ;
assign n3102 = (n46)*(n47) ;
assign n3103 = (n48)*((n46)*(n47)) ;
assign V321(2) = (~(((~((~((~(n617))*((~(n617))*(~(n647)))))*(~(n658))))*(n616))*(~((~(n616))*(~(n661))))))*(~(((n148)*(~(n616)))*((~(n616))*(~(n661)))));
assign V356 = ((~((n4994)*(n4997)))*(~((n5084)*(n5087))))*((n5214)*(n5216));
assign V357 = (~(n1218))*((n5990)*((n5992)*(~((n5540)*(n5544)))));
assign V373 = (n7)*(n8);
assign V375(0) = ~((n1286)*(((~((n53)*(n71)))*((~((n53)*(n163)))*(~((n53)*(n72)))))*(n1299)));
assign V377 = (n10)*(~((~(n9))*(~((n60)*((~(n59))*((n10)*(n65)))))));
assign V393(0) = ~((~((~(((~(n1389))*(~(n1395)))*((~(n1403))*(~(n1409)))))*(n6784)))*(n6831));
assign V398(0) = ~((~((~(((~(n1389))*(~(n1395)))*((~(n1403))*(~(n1409)))))*(n6784)))*(n7053));
assign V410(0) = ~(((~((~(n204))*(n205)))*(~((n204)*(n205))))*((~(n1308))*(~((n7118)*(~(n1474))))));
assign V423(0) = ~((((~(n1310))*(~((~(n489))*((~(n599))*(~(n629))))))*(n7016))*(n7019));
assign V432 = (~((~(((~(n1389))*(~(n1395)))*((~(n1403))*(~(n1409)))))*(n6784)))*(n7541);
assign V435(0) = ~((~(n1601))*(~(n1616)));
assign V500(0) = ~((~(n24))*(n151));
assign V508(0) = ~((n1622)*((~((n16)*(n559)))*(~(n1630))));
assign V511(0) = ~((~(n25))*(~((~(n21))*(n26))));
assign V512 = ((~((n251)*(~(n252))))*(~((~(n251))*(n252))))*((~((n249)*(~(n250))))*(~((~(n249))*(n250))));
assign V527 = ((((~(n21))*(~(n22)))*(~(n1308)))*(~(n1480)))*(~((n7746)*(n7745)));
assign V537 = ((~(n17))*(n508))*(~(n806));
assign V538 = ((~(n17))*(n508))*(~(n825));
assign V539 = ((~(n17))*(n508))*(~(n725));
assign V540 = ((~(n17))*(n508))*(~(n848));
assign V541 = ((~(n17))*(n508))*(~(n1679));
assign V542 = ((~(n17))*(n508))*(~(n1702));
assign V543 = ((~(n17))*(n508))*(~(n1725));
assign V544 = ((~(n17))*(n508))*(~(n1751));
assign V545 = ((~(n17))*(n508))*(~(n1777));
assign V546 = ((~(n17))*(n508))*(~(n1803));
assign V547 = ((~(n17))*(n508))*(~(n1830));
assign V548 = ((~(n17))*(n508))*(~(n1854));
assign V572(9) = ~((~((~(n1856))*((n1866)*(n1868))))*(~((~(n1871))*((~(n1866))*((~(n120))*(~(n1856)))))));
assign V572(8) = ~((~((~(n1383))*((n9048)*(n1866))))*(~((~(n1866))*((n9087)*(~(n1856))))));
assign V572(7) = ~((~(((n1866)*(~(n1364)))*(n9118)))*(~((~(n1856))*((n9181)*(~(n1866))))));
assign V572(6) = ~((~((~(n1920))*((n9304)*(n1866))))*(~((~(n1866))*((n9361)*(~(n1856))))));
assign V572(5) = ~((~((~(n1856))*((n1866)*(n1956))))*(~((~(n1871))*((~(n1866))*(n1964)))));
assign V572(4) = ~((~((~(n1856))*((n1866)*(n1991))))*(~((~(n1871))*((~(n1866))*((~(n1856))*(~(n1998)))))));
assign V572(3) = ~((~((~(n2030))*((n9924)*(n1866))))*(n2048));
assign V572(2) = ~((~((~(n2077))*((n10219)*(n1866))))*(n2095));
assign V572(1) = ~((~((~(n2124))*((n10517)*(n1866))))*(n2143));
assign V572(0) = ~((~((~(n667))*((n10663)*(n1866))))*((~((n1866)*(n10696)))*(~((n10750)*(~(n1866))))));
assign V585(0) = ~V34(0);
assign V587 = (~(n34))*(~((~((~(n70))*(~(n77))))*(~((~(n541))*((~(n484))*(~(n597)))))));
assign V591(0) = ~((~((~((~((~(n70))*(~(n77))))*(~((~(n541))*(n628)))))*((~(n34))*(n35))))*(~((~((~((~(n70))*(~(n77))))*(~((~(n541))*(n628)))))*((n34)*(~(n35))))));
assign V597(0) = ~((~((~((~((~(n70))*(~(n77))))*(~(n629))))*((n36)*(~((n34)*(n35))))))*(~((~((~((~(n70))*(~(n77))))*(~(n629))))*((~(n36))*((n34)*(n35))))));
assign V603(0) = ~((~((~((~(n489))*(~(n629))))*((n37)*(~((n36)*((n34)*(n35)))))))*(~((~((~(n489))*(~(n629))))*((~(n37))*((n36)*((n34)*(n35)))))));
assign V609(0) = ~((~((~((~(n489))*(~(n629))))*((n38)*(~((n37)*((n36)*(n1321)))))))*(~((~((~(n489))*(~(n629))))*((~(n38))*((n37)*((n36)*(n1321)))))));
assign V620 = (~(n2186))*((~((~(n1308))*(n2188)))*(~((~(n22))*((n1630)*((~(n1308))*(~(n1480)))))));
assign V621 = (n39)*((~((~(n26))*(n253)))*(~((n26)*(~(n253)))));
assign V630 = (~((n7589)*(~((~(n489))*(n1605)))))*(n7618);
assign V634(0) = (~((n43)*((~(n24))*(~((~(n24))*((n43)*(~(n44))))))))*(~((n42)*((n24)*(~((~(n24))*((n43)*(~(n44))))))));
assign V640(0) = ~((~(n24))*(~((~(n24))*((n43)*(~(n44))))));
assign V657 = ~V257(7);
assign V707 = (~(n57))*((~(n17))*((~(n55))*((~(n54))*(~(n56)))));
assign V763 = (~((~((n489)*((~(n68))*(~(n502)))))*((~(n508))*(~(n510)))))*(n3250);
assign V775 = ((n11480)*(n516))*(n2254);
assign V778 = (n53)*(n71);
assign V779 = (n72)*((n7)*(~(n8)));
assign V780 = (n53)*(n72);
assign V781 = (n72)*((n73)*(~((~(n70))*(~((~(n17))*((n5)*(~(n502))))))));
assign V782 = (n32)*((n7)*(~(n8)));
assign V783 = (n71)*(n74);
assign V784 = (n32)*(n74);
assign V787 = (n32)*(n53);
assign V789 = (n75)*((n53)*(~((~(n8))*((n44)*(n182)))));
assign V798(0) = ~((((~((n2276)*((~(n1421))*(~(n2298)))))*(n2307))*(~(n2338)))*(n11857));
assign V801 = ((~(n63))*((~(n61))*((n76)*((n20)*(~(n62))))))*(n502);
assign V802(0) = ~((~(n70))*(~(n77)));
assign V821(0) = ~((~((~(n80))*(~((~((~(n70))*(~(n77))))*((n57)*(n554))))))*(~((n29)*((~((~(n70))*(~(n77))))*((n57)*(n554))))));
assign V826(0) = ~((~((~(n81))*((~(n80))*(~((~(n489))*((n57)*(n554)))))))*((~((n80)*((n81)*(~((~(n489))*((n57)*(n554)))))))*(~((n30)*((~(n489))*((n57)*(n554)))))));
assign V966 = (n151)*((n2254)*(~((~((~((~(n70))*(~(n77))))*(~(n2338))))*(n12005))));
assign V986 = (n151)*((n2254)*(~((~(n2365))*((~((n15)*(~(n537))))*(~(n2369))))));
assign V1213(11) = ~((~((n616)*((~((~(n616))*(~(n661))))*(~((~(n1842))*(~(n1848)))))))*(~(((n136)*(~(n616)))*((~(n616))*(~(n661))))));
assign V1213(10) = ~((~((n616)*((~((~(n616))*(~(n661))))*(~((~(n1818))*(~(n1824)))))))*(~(((n137)*(~(n616)))*((~(n616))*(~(n661))))));
assign V1213(9) = ~((~(((~(n1798))*(n616))*(~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))))*(~((~(n616))*((n138)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))));
assign V1213(8) = ~((~(((~(n1772))*(n616))*(~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))))*(~((~(n616))*((n131)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))));
assign V1213(7) = ~((~(((~(n1746))*(n616))*(~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))))*(~((~(n616))*((n132)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))));
assign V1213(6) = ~((~(((~((~((~(n617))*((~(n617))*(~(n1715)))))*(~((n617)*((n617)*(n652))))))*(n616))*(~((~(n616))*(~(n661))))))*(~(((n133)*(~(n616)))*((~(n616))*(~(n661))))));
assign V1213(5) = ~((~(((~((~((~(n617))*((~(n617))*(~(n1692)))))*(~((n617)*((n617)*(~(n652)))))))*(n616))*(~((~(n616))*(~(n661))))))*(~(((n134)*(~(n616)))*((~(n616))*(~(n661))))));
assign V1213(4) = ~((~((((~((n516)*(n537)))*(~((~(n616))*(~(n661)))))*(n616))*(~(n1672))))*(~(((n135)*(~(n616)))*((~(n616))*(~(n661))))));
assign V1213(3) = ~((~((n616)*((~((~(n616))*(~(n661))))*(n843))))*(~(((n4)*(~(n616)))*((~(n616))*(~(n661))))));
assign V1213(2) = ~((~((n616)*((~((~(n616))*(~(n661))))*(n720))))*(~(((n3)*(~(n616)))*((~(n616))*(~(n661))))));
assign V1213(1) = ~((~((n616)*((~((~(n616))*(~(n661))))*(n820))))*(~(((n2)*(~(n616)))*((~(n616))*(~(n661))))));
assign V1213(0) = ~((~((n616)*((~((~(n616))*(~(n661))))*(n801))))*(~(((n1)*(~(n616)))*((~(n616))*(~(n661))))));
assign V1243(9) = ~((~((n616)*((~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))*(~(n1340)))))*(~((~(n616))*((n139)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))));
assign V1243(8) = ~((~((n616)*((~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))*(~(n1378)))))*(~((~(n616))*((n140)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))));
assign V1243(7) = ~((~((n616)*((~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))*(~(n1359)))))*(~((~(n616))*((n141)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))));
assign V1243(6) = ~((~((n616)*((~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))*(~(n1915)))))*(~((~(n616))*((n142)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))));
assign V1243(5) = ~((~((n616)*((~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))*(~(n1949)))))*(~((~(n616))*((n143)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))));
assign V1243(4) = ~((~((n616)*((~((~(n616))*(~((n164)*(~((~(n595))*(~(n597))))))))*(~(n1984)))))*(~((~(n616))*((n144)*((~(n616))*(~((n164)*(~((~(n595))*(~(n597)))))))))));
assign V1243(3) = ~((~((n616)*((~((~(n616))*(~(n661))))*(~((~(n2018))*(~(n2024)))))))*(~(((n145)*(~(n616)))*((~(n616))*(~(n661))))));
assign V1243(2) = ~((~((n616)*((~((~(n616))*(~(n661))))*(~((~(n2065))*(~(n2071)))))))*(~(((n146)*(~(n616)))*((~(n616))*(~(n661))))));
assign V1243(1) = ~((~((n616)*((~((~(n616))*(~(n661))))*(~((~(n2112))*(~(n2118)))))))*(~(((n147)*(~(n616)))*((~(n616))*(~(n661))))));
assign V1243(0) = ~((~(((~((~((~(n617))*((~(n617))*(~(n647)))))*(~(n658))))*(n616))*(~((~(n616))*(~(n661))))))*(~(((n148)*(~(n616)))*((~(n616))*(~(n661))))));
assign V1256 = (n149)*((n7)*(~(n8)));
assign V1257 = (n12198)*((~((n166)*(~(((n12134)*(n587))*(n1430)))))*(~((~(n166))*(n1535))));
assign V1258 = (n53)*(n149);
assign V1259 = (n53)*(n150);
assign V1260 = (n74)*(n150);
assign V1261 = (~(n15))*((n74)*(n150));
assign V1262 = (n75)*((n7)*(~(n8)));
assign V1263 = (n53)*(n75);
assign V1264 = (n73)*(n75);
assign V1265 = (n70)*((n73)*(n75));
assign V1266 = (n74)*(n75);
assign V1267 = (n74)*(n149);
assign V1274(0) = ~((~(((n15)*((n151)*(n2254)))*(n559)))*(~((n2254)*((n12333)*(n12337)))));
assign V1281(0) = ~((~(((~((~((n12414)*(~(n2419))))*(n12486)))*(~(n2428)))*(n12496)))*(~((~((~((~((n12414)*(~(n2419))))*(n12486)))*(~(n2428))))*((~((~((~((n12414)*(~(n2419))))*(n12486)))*(~(n2428))))*(~(n2439))))));
assign V1297(4) = ~((~(((n153)*(~(n2428)))*((n151)*(~((n5)*(n2279))))))*(~((n2428)*((n64)*(n2428)))));
assign V1297(3) = ~((~(((n154)*(~(n2428)))*((n151)*(~((n5)*(n2279))))))*(~((n2428)*((n63)*(n2428)))));
assign V1297(2) = ~((~(((n155)*(~(n2428)))*((n151)*(~((n5)*(n2279))))))*(~((n2428)*((n62)*(n2428)))));
assign V1297(1) = ~((~(((n156)*(~(n2428)))*((n151)*(~((n5)*(n2279))))))*(~((n2428)*((n61)*(n2428)))));
assign V1297(0) = ~((~(((n157)*(~(n2428)))*((n151)*(~((n5)*(n2279))))))*(~((n2428)*((n76)*(n2428)))));
assign V1365 = (((~((n28)*(n1569)))*(~((~(n28))*(n1569))))*((~(n1535))*((n151)*(n2254))))*(n12619);
assign V1375 = ~V268(5);
assign V1378 = ((n32)*((n7)*(~(n8))))*((~((~(n70))*(~(n77))))*(~(n628)));
assign V1380 = ((n32)*((n7)*(~(n8))))*(~((n12776)*(~(n1865))));
assign V1382 = ((n7)*(~(n8)))*((n32)*(~((~(n595))*(~((~(n489))*(~(n1539)))))));
assign V1384 = (((n7)*(~(n8)))*(~((~(n1529))*(~((~(n1538))*(~(n1541)))))))*(n12818);
assign V1386 = ((n7)*(~(n8)))*((n32)*((~((~(n193))*(n536)))*(~(n2508))));
assign V1387 = (n53)*(n163);
assign V1392(0) = ~((~(((n151)*(n2254))*((n12891)*(n516))))*(~(((n151)*(n2254))*(n12949))));
assign V1423 = (n31)*(n53);
assign V1426 = (n31)*((n7)*(~(n8)));
assign V1428 = (n31)*(n74);
assign V1429 = (n31)*(n73);
assign V1431 = ((n31)*(n53))*(~((~(n8))*(n167)));
assign V1432 = (n151)*((n19)*(n2254));
assign V1439(0) = ~((~((~(n28))*((n30)*(n494))))*(~((n151)*((n168)*(~(n597))))));
assign V1440(0) = ~((n151)*(~((n169)*(~((n168)*((~(n17))*(n508)))))));
assign V1451(0) = ~((~((n85)*((n151)*((~((~((~(n193))*(n536)))*(~(n2508))))*(~(n2535))))))*(~((~(n85))*((n151)*(~((~((~((~(n193))*(n536)))*(~(n2508))))*(~(n2535))))))));
assign V1459(0) = ~((~((n151)*((n170)*((~((~(n85))*((~(n537))*(~(n2508)))))*(~((n85)*(n2535)))))))*(~((n151)*((~(n170))*(~((~((~(n85))*((~(n537))*(~(n2508)))))*(~((n85)*(n2535)))))))));
assign V1467(0) = ~((~((n151)*((n171)*((~((~(n170))*((~(n85))*(n2509))))*(~((n170)*((n85)*(n2535))))))))*(~((n151)*((~(n171))*(~((~((~(n170))*((~(n85))*(n2509))))*(~((n170)*((n85)*(n2535))))))))));
assign V1470 = (n172)*((n2254)*((n151)*(~(n1580))));
assign V1480(0) = ~((~((~(n554))*(~(n1472))))*((~((~(n1529))*(~((~(n1538))*(~(n1541))))))*(~(((n554)*(~(n1472)))*(~(n489))))));
assign V1481(0) = ~V214(0);
assign V1492(0) = ~((~((~(n22))*(n175)))*(~((n2246)*(n2571))));
assign V1495(0) = ~V175(0);
assign V1512(3) = ~((~((n2249)*(~((n13312)*(n2249)))))*(~(((n13312)*(n2249))*(~((~((n5540)*(n5544)))*((n13382)*(n13385)))))));
assign V1512(2) = ~((~((~(n2591))*(~((n13402)*(n2249)))))*(~((n2591)*(~((n2605)*((n13453)*(n13455)))))));
assign V1512(1) = ~((~((~(n2591))*(~((n2249)*(n2261)))))*(~((n2591)*(~((n2605)*((n13513)*(n13515)))))));
assign V1536(0) = ~((n13312)*(n2249));
assign V1537 = (n151)*((n173)*(n2254));
assign V1539 = (n151)*((n2254)*(~((~(n174))*(~(n180)))));
assign V1552(1) = ~((~((((~(n110))*(~((~(n489))*(~(n1539)))))*(n595))*(n489)))*(~(((~(n489))*(~(n1539)))*((~(n1345))*(~((n489)*(n595)))))));
assign V1552(0) = ~((~(n2641))*(~(((~(n489))*(~(n1539)))*((~(n1383))*(~((n489)*(n595)))))));
assign V1613(0) = (~((~(n2696))*(n2781)))*(~((n2696)*(~(n2781))));
assign V1613(1) = (~((~((~((~((~((~(n2789))*(n2794)))*(~((n2789)*(~(n2794))))))*((~((~(n2804))*(n2811)))*(~((n2804)*(~(n2811)))))))*(~(((~((~(n2789))*(n2794)))*(~((n2789)*(~(n2794)))))*(~((~((~(n2804))*(n2811)))*(~((n2804)*(~(n2811))))))))))*((~((~(n2834))*(n2851)))*(~((n2834)*(~(n2851)))))))*(~(((~((~((~((~(n2789))*(n2794)))*(~((n2789)*(~(n2794))))))*((~((~(n2804))*(n2811)))*(~((n2804)*(~(n2811)))))))*(~(((~((~(n2789))*(n2794)))*(~((n2789)*(~(n2794)))))*(~((~((~(n2804))*(n2811)))*(~((n2804)*(~(n2811)))))))))*(~((~((~(n2834))*(n2851)))*(~((n2834)*(~(n2851))))))));
assign V1620(0) = ~(((~(n488))*(~((n17)*(~(n2249)))))*(n15300));
assign V1629(0) = ~((~((~((n1535)*(~((~(n1529))*(~((~(n1538))*(~(n1541))))))))*(n2864)))*(n2870));
assign V1645(0) = ~((~((~((~((n7223)*(n1546)))*(n7294)))*(~((n7380)*(n7378)))))*(n2873));
assign V1652(0) = ~((~(n79))*((n189)*((~(n1605))*((~(n14))*((~(n6))*(n537))))));
assign V1669 = (~((n489)*(n2880)))*((~(((n2249)*(n2298))*(n15570)))*(n2904));
assign V1671(0) = ~V205(0);
assign V1679(0) = ~((n536)*(~((n15443)*(n193))));
assign V1693(0) = ~((~(((~(n2910))*(~((~((n12414)*(~(n2419))))*(n15681))))*(n15693)))*(~((~((~(n2910))*(~((~((n12414)*(~(n2419))))*(n15681)))))*((~(n2439))*(~((~(n2910))*(~((~((n12414)*(~(n2419))))*(n15681)))))))));
assign V1709(4) = ~((~(((n195)*((n151)*(~((n5)*(n2282)))))*(~(n2910))))*(~((n2910)*((n64)*(n2910)))));
assign V1709(3) = ~((~(((n196)*((n151)*(~((n5)*(n2282)))))*(~(n2910))))*(~((n2910)*((n63)*(n2910)))));
assign V1709(2) = ~((~(((n197)*((n151)*(~((n5)*(n2282)))))*(~(n2910))))*(~((n2910)*((n62)*(n2910)))));
assign V1709(1) = ~((~(((n198)*((n151)*(~((n5)*(n2282)))))*(~(n2910))))*(~((n2910)*((n61)*(n2910)))));
assign V1709(0) = ~((~(((n199)*((n151)*(~((n5)*(n2282)))))*(~(n2910))))*(~((n2910)*((n76)*(n2910)))));
assign V1717(0) = ~((~((n2254)*(n15834)))*(~((~(n489))*(~(n2960)))));
assign V1719 = (~(n178))*((n200)*(~((n65)*((n59)*(~(n60))))));
assign V1726(0) = ~((~((n628)*((n151)*(n201))))*(~((n2591)*((~(n629))*(n1859)))));
assign V1736 = (~(n79))*((n489)*(((~(n541))*(~((n202)*(~(n628)))))*(n2880)));
assign V1741(0) = ~(((~((n79)*(n1308)))*(~(n2240)))*((n11541)*(~((~(n1308))*(n2235)))));
assign V1745(0) = ~((~(n508))*((n6)*((n203)*(~((n28)*((n30)*(n499)))))));
assign V1757(0) = ~((~((~(n204))*(n205)))*(~(n1471)));
assign V1758(0) = ~((~((~(n204))*(n205)))*(~((n204)*(~(n205)))));
assign V1759(0) = ~((~((n151)*((n206)*(~((n5)*((n28)*(n832)))))))*(n2981));
assign V1760(0) = ~V101(0);
assign V1771(1) = ~((~(((n28)*(n549))*((~(n67))*((n28)*(n549)))))*(~((~((n28)*(n549)))*((~(n244))*(~((n28)*(n549)))))));
assign V1771(0) = ~((~(((n28)*(n549))*((~(n66))*((n28)*(n549)))))*(~((~((n28)*(n549)))*((~(n245))*(~((n28)*(n549)))))));
assign V1781(1) = ~((~((~((n28)*(n549)))*((~((n28)*(n549)))*(n1854))))*(~(((n28)*(n549))*((~(n248))*((n28)*(n549))))));
assign V1781(0) = ~((~((~((n28)*(n549)))*((~((n28)*(n549)))*(n1830))))*(~(((n28)*(n549))*((~(n247))*((n28)*(n549))))));
assign V1829(9) = ~((~((n23)*((n23)*(n1345))))*(~((~(n23))*((~(n23))*(n667)))));
assign V1829(8) = ~((~((n23)*((n23)*(n1383))))*(~((~(n23))*((~(n23))*(n1854)))));
assign V1829(7) = ~((~((n23)*((n23)*(n1364))))*(~((~(n23))*((~(n23))*(n1830)))));
assign V1829(6) = ~((~((n23)*((n23)*(n1920))))*(~((~(n23))*((~(n23))*(n1803)))));
assign V1829(5) = ~((~((n23)*((n23)*(n1954))))*(~((~(n23))*((~(n23))*(n1777)))));
assign V1829(4) = ~((~((n23)*((n23)*(n1989))))*(~((~(n23))*((~(n23))*(n1751)))));
assign V1829(3) = ~((~((n23)*((n23)*(n2030))))*(~((~(n23))*((~(n23))*(n1725)))));
assign V1829(2) = ~((~((n23)*((n23)*(n2077))))*(~((~(n23))*((~(n23))*(n1702)))));
assign V1829(1) = ~((~((n23)*((n23)*(n2124))))*(~((~(n23))*((~(n23))*(n1679)))));
assign V1829(0) = ~((~((~(n23))*((~(n23))*(n667))))*(~((n23)*((n23)*(n725)))));
assign V1832 = (n151)*(~((~(n2535))*(~((n192)*(~((~(n2508))*((n193)*(~((n15443)*(n193))))))))));
assign V1833(0) = ~V261(0);
assign V1863(0) = ~V301(0);
assign V1864(0) = ~V302(0);
assign V1896(0) = ~(((~(n1471))*(~((~(n1529))*(~((~(n1538))*(~(n1541)))))))*(~((n212)*(~(n3056)))));
assign V1897(0) = ~((~((n597)*((~(n1529))*(~((~(n1538))*(~(n1541)))))))*(~((n213)*(~(n3056)))));
assign V1898(0) = ~((~((n508)*(n2230)))*(~((n214)*(~((n5)*(n2322))))));
assign V1899(0) = ~((~((n510)*(n2230)))*(~((n215)*(~((n5)*(n2322))))));
assign V1900(0) = ~((~((~(n204))*(n205)))*(~((n216)*(~((n5)*(n2322))))));
assign V1901(0) = ~((~((n204)*(~(n205))))*(~((n217)*(~((n5)*((n28)*(n832)))))));
assign V1921(5) = ~((~((n218)*((n13795)*(n2287))))*(n2670));
assign V1921(4) = ~((n2680)*(n2689));
assign V1921(3) = ~((n2705)*(n2714));
assign V1921(2) = ~((n2724)*(n2733));
assign V1921(1) = ~((n2746)*(n2755));
assign V1921(0) = ~((n2765)*(n2774));
assign V1953(1) = (~((n28)*(n832)))*((~((~(n28))*(n549)))*((n230)*((~(n28))*(n1532))));
assign V1953(7) = ~((~((~((n28)*(n832)))*((~((~(n28))*(n549)))*((n224)*((~(n28))*(n1532))))))*(~((~((n28)*(n832)))*(((~(n28))*(n549))*((n232)*(~((~(n28))*(n1532))))))));
assign V1953(6) = ~((~((~((n28)*(n832)))*((~((~(n28))*(n549)))*((n225)*((~(n28))*(n1532))))))*(~((~((n28)*(n832)))*(((~(n28))*(n549))*((n233)*(~((~(n28))*(n1532))))))));
assign V1953(5) = ~((~((~((n28)*(n832)))*((~((~(n28))*(n549)))*((n226)*((~(n28))*(n1532))))))*(~((~((n28)*(n832)))*(((~(n28))*(n549))*((n234)*(~((~(n28))*(n1532))))))));
assign V1953(4) = ~((~((~((n28)*(n832)))*((~((~(n28))*(n549)))*((n227)*((~(n28))*(n1532))))))*(~((~((n28)*(n832)))*(((~(n28))*(n549))*((n235)*(~((~(n28))*(n1532))))))));
assign V1953(3) = ~((~((~((n28)*(n832)))*((~((~(n28))*(n549)))*((n228)*((~(n28))*(n1532))))))*(~((~((n28)*(n832)))*(((~(n28))*(n549))*((n236)*(~((~(n28))*(n1532))))))));
assign V1953(2) = ~((~((~((n28)*(n832)))*((~((~(n28))*(n549)))*((n229)*((~(n28))*(n1532))))))*(~((~((n28)*(n832)))*(((~(n28))*(n549))*((n237)*(~((~(n28))*(n1532))))))));
assign V1953(0) = ~((~((~((n28)*(n832)))*((~((~(n28))*(n549)))*((n231)*((~(n28))*(n1532))))))*(~(((n28)*(n832))*((~((~(n28))*(n549)))*((n217)*(~((~(n28))*(n1532))))))));
assign V1960(1) = ~((~((n238)*(((~(n1566))*(~((n28)*(n1569))))*((~(n28))*(n549)))))*(~((n240)*((~((~(n1566))*(~((n28)*(n1569)))))*(~((~(n28))*(n549)))))));
assign V1960(0) = ~((~((n239)*(((~(n1566))*(~((n28)*(n1569))))*((~(n28))*(n549)))))*(~((n241)*((~((~(n1566))*(~((n28)*(n1569)))))*(~((~(n28))*(n549)))))));
assign V1968(0) = ~((~((~((n5)*((~(n28))*(n549))))*(n16040)))*(~((~(n243))*(n16087))));
assign V1992(1) = ~((~((~((~(n1861))*(~((~(n489))*(~(n628))))))*((n1861)*((~(n244))*(~((~(n489))*(~(n628))))))))*(~((~((n1861)*(~((~(n489))*(~(n628))))))*((~((~(n489))*(~(n628))))*((n244)*(~(n1861)))))));
assign V1992(0) = ~((~((~((~(n1861))*(~((~(n489))*(~(n628))))))*((n1861)*((~((~(n489))*(~(n628))))*(~((~((n244)*(~(n245))))*(~((~(n244))*(n245)))))))))*(~((~((n1861)*(~((~(n489))*(~(n628))))))*((~((~(n489))*(~(n628))))*((n245)*(~(n1861)))))));
assign V650 = ~((~((n130)*(~((n52)*((n51)*((n50)*((n49)*(n3103))))))))*(~((~(n130))*((n52)*((n51)*((n50)*((n49)*(n3103))))))));
assign V651 = ~((~((n49)*(~((n52)*((n51)*((n50)*((n48)*(n3102))))))))*(~((~(n49))*((n52)*((n51)*((n50)*((n48)*(n3102))))))));
assign V652 = ~((~((n50)*(~((n52)*((n51)*((n48)*((n46)*(n47))))))))*(~((~(n50))*((n52)*((n51)*((n48)*((n46)*(n47))))))));
assign V653 = ~((~((n48)*(~((n52)*((n51)*((n46)*(n47)))))))*(~((~(n48))*((n52)*((n51)*((n46)*(n47)))))));
assign V654 = ~((~((n51)*(~((n52)*((n46)*(n47))))))*(~((~(n51))*((n52)*((n46)*(n47))))));
assign V655 = ~((~((n47)*(~((n46)*(n52)))))*(~((~(n47))*((n46)*(n52)))));
assign V656 = ~((~((~(n46))*(n52)))*(~((n46)*(~(n52)))));
assign V1370 = ~((~((n207)*(~((n162)*((n161)*((n160)*((n158)*(n159))))))))*(~((~(n207))*((n162)*((n161)*((n160)*((n158)*(n159))))))));
assign V1371 = ~((~((n160)*(~((n162)*((n161)*((n158)*(n159)))))))*(~((~(n160))*((n162)*((n161)*((n158)*(n159)))))));
assign V1372 = ~((~((n161)*(~((n162)*((n158)*(n159))))))*(~((~(n161))*((n162)*((n158)*(n159))))));
assign V1373 = ~((~((n159)*(~((n158)*(n162)))))*(~((~(n159))*((n158)*(n162)))));
assign V1374 = ~((~((~(n158))*(n162)))*(~((n158)*(~(n162)))));
endmodule

